module Sobol_to_INT32(
    input             clk,
    input             rst_n, 
    input             start,
    output reg [31:0] res
);
// ================== parameter =========================
parameter IDLE = 1'b0;
parameter COMP = 1'b1;
// DVA31, DVA30 , ......, DVA1, DVA0
parameter [32*32-1:0] DVA = {
    32'b00000000000000000000000111110011,
    32'b00000000000000000000001100110010,
    32'b00000000000000000000011011000100,
    32'b00000000000000000000110110001000,
    32'b00000000000000000001101111010000,
    32'b00000000000000000011011101100000,
    32'b00000000000000000110111101000000,
    32'b00000000000000001101111110000000,
    32'b00000000000000000100110100000000,
    32'b00000000000000000100111000000000,
    32'b00000000000000000011110000000000,
    32'b00000000000000000111100000000000,
    32'b00000000000000000011000000000000,
    32'b00000000000000001010000000000000,
    32'b00000000000000001100000000000000,
    32'b00000000000000001000000000000000,
    32'b00000001111100110000000000000000,
    32'b00000011001100100000000000000000,
    32'b00000110110001000000000000000000,
    32'b00001101100010000000000000000000,
    32'b00011011110100000000000000000000,
    32'b00110111011000000000000000000000,
    32'b01101111010000000000000000000000,
    32'b11011111100000000000000000000000,
    32'b01001101000000000000000000000000,
    32'b01001110000000000000000000000000,
    32'b00111100000000000000000000000000,
    32'b01111000000000000000000000000000,
    32'b00110000000000000000000000000000,
    32'b10100000000000000000000000000000,
    32'b11000000000000000000000000000000,
    32'b10000000000000000000000000000000
};


// ================== reg and wire ======================
// reg   [31:0] res0, res1, res2, res3;
wire  [31:0] res_w;

reg          state, state_ns;

reg   [31:0] counter;
reg   [4:0] LSZ;

integer i;

// ================== wire assignments ==================
assign res_w = res ^ DVA[32*(LSZ+1)-1 -: 32];

// ================== Combinational =====================
// state
always @(*) begin
    state_ns = state;
    case (state_ns)
        IDLE: begin
            if (start) state_ns = COMP;
        end 
        COMP: begin
            
        end
        default: begin
            
        end
    endcase
end
// counter 
always @(*) begin
    for (i=0; i < 32; i = i+1) begin
        if (counter[31 - i] == 0) LSZ = 31 - i;
    end
end


// ================== sequential ========================
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        res     <= 32'b0;
        counter <= 32'b0;
        state   <= IDLE;
    end
    else begin
        state <= state_ns;
        if (state == COMP) begin
            res     <= res_w;
            counter <= counter + 32'b1;
        end
        else begin
            res     <= 32'b0;
            counter <= 32'b0;
        end
    end
end

endmodule