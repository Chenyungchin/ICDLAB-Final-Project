* SPICE NETLIST
***************************************

.SUBCKT L POS NEG SUB
.ENDS
***************************************
.SUBCKT YA2GSD O E2 E8 E4 I SR E
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=0
X0 1 2 2 2 5 3 4 YA2GSD $T=0 0 0 0 $X=2850 $Y=0
.ENDS
***************************************
.SUBCKT XMD I SMT PU PD O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4
** N=4 EP=4 IP=6 FDC=0
X0 1 2 2 2 3 XMD $T=0 0 0 0 $X=2850 $Y=0
.ENDS
***************************************
.SUBCKT ICV_3 1 2 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 30 31 32
+ 33 34 49
** N=69 EP=23 IP=48 FDC=0
X0 11 1 1 1 34 XMD $T=243040 1350160 0 180 $X=183270 $Y=1210660
X1 12 1 1 1 21 XMD $T=345960 1350160 0 180 $X=286190 $Y=1210660
X2 13 14 14 14 22 XMD $T=448880 1350160 0 180 $X=389110 $Y=1210660
X3 15 2 2 2 23 XMD $T=551800 1350160 0 180 $X=492030 $Y=1210660
X4 16 9 9 9 30 XMD $T=860560 1350160 0 180 $X=800790 $Y=1210660
X5 17 9 9 9 31 XMD $T=963480 1350160 0 180 $X=903710 $Y=1210660
X6 18 10 10 10 32 XMD $T=1066400 1350160 0 180 $X=1006630 $Y=1210660
X7 19 20 20 20 33 XMD $T=1169320 1350160 0 180 $X=1109550 $Y=1210660
.ENDS
***************************************
.SUBCKT INV1S I VCC O GND
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF1S I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DELB I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DELA I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT QDFFRBN D CK RB VCC GND Q
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=0
X0 1 2 3 4 DELB $T=0 0 0 0 $X=0 $Y=-380
X1 5 2 3 6 DELB $T=4960 0 0 0 $X=4960 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=0
X0 1 2 3 4 DELB $T=0 0 0 0 $X=0 $Y=-380
X1 5 2 3 6 DELA $T=4960 0 0 0 $X=4960 $Y=-380
.ENDS
***************************************
.SUBCKT MUX2 B S VCC GND O A
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22S A1 B1 O B2 GND A2 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN4S I1 I2 I4 I3 VCC GND O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF1 I VCC GND O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF1CK I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV2 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF2 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND3 I3 GND I2 O VCC I1
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND2S I1 O I2 VCC GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MOAI1S B1 B2 GND A1 A2 O VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR2 I1 VCC O I2 GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV12CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2 I2 I1 VCC GND O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA22 A1 A2 B1 B2 VCC GND O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN2 I1 I2 GND VCC O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR3 I1 VCC I2 I3 O GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2B1S I1 B1 GND O VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 247 248 249 250 251 252 253 254 255 256 257 259 260 261 262 263
+ 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283
+ 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 301 302 303 304
+ 305 306 307 309 310 311 312 313 314 315 316 317 319 320 321 322 323 324 325 326
+ 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342 343 344 345 346
+ 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362 363 364 365 366
+ 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382 383 384 385 386
+ 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406
+ 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426
+ 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446
+ 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466
+ 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486
+ 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506
+ 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526
+ 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546
+ 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566
+ 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586
+ 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606
+ 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626
+ 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646
+ 647 648 649 650 651 652 653 667 681
** N=1339 EP=649 IP=5627 FDC=0
X0 652 1338 1338 1338 667 651 653 YA2GSD $T=1349740 1096780 0 90 $X=1210240 $Y=1099630
X1 10 2 685 1 INV1S $T=306280 1092120 0 180 $X=305040 $Y=1086700
X2 690 2 695 1 INV1S $T=316820 1102200 1 0 $X=316820 $Y=1096780
X3 17 2 707 1 INV1S $T=344720 1102200 1 0 $X=344720 $Y=1096780
X4 710 2 712 1 INV1S $T=349060 1102200 0 0 $X=349060 $Y=1101820
X5 21 2 713 1 INV1S $T=352780 1092120 1 0 $X=352780 $Y=1086700
X6 714 2 709 1 INV1S $T=356500 1112280 0 180 $X=355260 $Y=1106860
X7 694 2 31 1 INV1S $T=367040 1092120 0 0 $X=367040 $Y=1091740
X8 31 2 722 1 INV1S $T=372000 1092120 0 0 $X=372000 $Y=1091740
X9 52 2 40 1 INV1S $T=410440 1092120 1 0 $X=410440 $Y=1086700
X10 52 2 747 1 INV1S $T=411680 1092120 1 0 $X=411680 $Y=1086700
X11 771 2 775 1 INV1S $T=455080 1102200 0 0 $X=455080 $Y=1101820
X12 88 2 76 1 INV1S $T=456940 1092120 0 180 $X=455700 $Y=1086700
X13 30 2 88 1 INV1S $T=455700 1092120 0 0 $X=455700 $Y=1091740
X14 774 2 777 1 INV1S $T=456940 1102200 0 0 $X=456940 $Y=1101820
X15 88 2 767 1 INV1S $T=458180 1092120 1 0 $X=458180 $Y=1086700
X16 781 2 784 1 INV1S $T=464380 1092120 1 0 $X=464380 $Y=1086700
X17 776 2 792 1 INV1S $T=473680 1092120 1 0 $X=473680 $Y=1086700
X18 801 2 132 1 INV1S $T=487320 1112280 1 0 $X=487320 $Y=1106860
X19 804 2 137 1 INV1S $T=493520 1092120 0 180 $X=492280 $Y=1086700
X20 807 2 138 1 INV1S $T=494760 1102200 0 0 $X=494760 $Y=1101820
X21 809 2 141 1 INV1S $T=500340 1092120 0 180 $X=499100 $Y=1086700
X22 811 2 118 1 INV1S $T=500960 1102200 1 180 $X=499720 $Y=1101820
X23 811 2 789 1 INV1S $T=500960 1102200 0 0 $X=500960 $Y=1101820
X24 811 2 153 1 INV1S $T=511500 1102200 0 0 $X=511500 $Y=1101820
X25 170 2 811 1 INV1S $T=529480 1092120 1 180 $X=528240 $Y=1091740
X26 847 2 836 1 INV1S $T=554900 1112280 0 180 $X=553660 $Y=1106860
X27 135 2 847 1 INV1S $T=555520 1112280 1 0 $X=555520 $Y=1106860
X28 207 2 822 1 INV1S $T=567300 1102200 1 0 $X=567300 $Y=1096780
X29 847 2 867 1 INV1S $T=577840 1112280 1 0 $X=577840 $Y=1106860
X30 205 2 876 1 INV1S $T=590860 1112280 1 0 $X=590860 $Y=1106860
X31 876 2 225 1 INV1S $T=592720 1102200 0 0 $X=592720 $Y=1101820
X32 189 2 233 1 INV1S $T=597680 1092120 1 0 $X=597680 $Y=1086700
X33 876 2 869 1 INV1S $T=599540 1112280 0 180 $X=598300 $Y=1106860
X34 233 2 885 1 INV1S $T=603260 1092120 0 0 $X=603260 $Y=1091740
X35 883 2 888 1 INV1S $T=604500 1112280 1 0 $X=604500 $Y=1106860
X36 874 2 892 1 INV1S $T=610080 1092120 0 0 $X=610080 $Y=1091740
X37 895 2 897 1 INV1S $T=611940 1112280 0 0 $X=611940 $Y=1111900
X38 903 2 906 1 INV1S $T=623720 1102200 1 180 $X=622480 $Y=1101820
X39 866 2 905 1 INV1S $T=624340 1092120 1 180 $X=623100 $Y=1091740
X40 219 2 263 1 INV1S $T=639220 1092120 1 0 $X=639220 $Y=1086700
X41 924 2 925 1 INV1S $T=642940 1102200 1 0 $X=642940 $Y=1096780
X42 920 2 928 1 INV1S $T=645420 1092120 1 0 $X=645420 $Y=1086700
X43 919 2 932 1 INV1S $T=647900 1112280 1 0 $X=647900 $Y=1106860
X44 940 2 938 1 INV1S $T=657200 1112280 0 180 $X=655960 $Y=1106860
X45 942 2 945 1 INV1S $T=663400 1102200 0 180 $X=662160 $Y=1096780
X46 950 2 952 1 INV1S $T=673320 1102200 1 180 $X=672080 $Y=1101820
X47 958 2 962 1 INV1S $T=681380 1112280 1 0 $X=681380 $Y=1106860
X48 960 2 929 1 INV1S $T=683860 1092120 0 0 $X=683860 $Y=1091740
X49 294 2 960 1 INV1S $T=685720 1092120 0 0 $X=685720 $Y=1091740
X50 301 2 971 1 INV1S $T=697500 1102200 0 180 $X=696260 $Y=1096780
X51 972 2 977 1 INV1S $T=699980 1122360 1 0 $X=699980 $Y=1116940
X52 985 2 987 1 INV1S $T=712380 1122360 1 0 $X=712380 $Y=1116940
X53 301 2 992 1 INV1S $T=713000 1092120 0 0 $X=713000 $Y=1091740
X54 996 2 994 1 INV1S $T=716100 1112280 1 180 $X=714860 $Y=1111900
X55 1003 2 1004 1 INV1S $T=723540 1112280 0 0 $X=723540 $Y=1111900
X56 993 2 1008 1 INV1S $T=726020 1092120 0 0 $X=726020 $Y=1091740
X57 1014 2 1016 1 INV1S $T=730980 1122360 1 0 $X=730980 $Y=1116940
X58 1009 2 314 1 INV1S $T=734700 1092120 1 180 $X=733460 $Y=1091740
X59 338 2 1060 1 INV1S $T=778100 1102200 1 0 $X=778100 $Y=1096780
X60 1060 2 334 1 INV1S $T=779340 1102200 1 0 $X=779340 $Y=1096780
X61 1060 2 1045 1 INV1S $T=780580 1102200 1 180 $X=779340 $Y=1101820
X62 1060 2 1073 1 INV1S $T=796700 1112280 0 180 $X=795460 $Y=1106860
X63 1060 2 351 1 INV1S $T=797940 1092120 1 180 $X=796700 $Y=1091740
X64 395 2 1142 1 INV1S $T=865520 1092120 1 180 $X=864280 $Y=1091740
X65 395 2 396 1 INV1S $T=865520 1092120 1 0 $X=865520 $Y=1086700
X66 396 2 409 1 INV1S $T=886600 1092120 1 0 $X=886600 $Y=1086700
X67 409 2 1165 1 INV1S $T=895280 1092120 0 0 $X=895280 $Y=1091740
X68 464 2 1214 1 INV1S $T=953560 1092120 1 0 $X=953560 $Y=1086700
X69 1214 2 1218 1 INV1S $T=956040 1092120 0 0 $X=956040 $Y=1091740
X70 525 2 373 1 INV1S $T=1020520 1122360 1 180 $X=1019280 $Y=1121980
X71 525 2 538 1 INV1S $T=1035400 1122360 0 0 $X=1035400 $Y=1121980
X72 551 2 1290 1 INV1S $T=1045320 1102200 1 0 $X=1045320 $Y=1096780
X73 1290 2 1292 1 INV1S $T=1049040 1102200 1 0 $X=1049040 $Y=1096780
X74 569 2 1309 1 INV1S $T=1071980 1092120 0 0 $X=1071980 $Y=1091740
X75 1309 2 583 1 INV1S $T=1074460 1092120 0 0 $X=1074460 $Y=1091740
X76 1309 2 1311 1 INV1S $T=1076940 1092120 0 0 $X=1076940 $Y=1091740
X77 525 2 1338 1 INV1S $T=1127780 1112280 0 0 $X=1127780 $Y=1111900
X78 707 1 2 19 BUF1S $T=344100 1102200 1 180 $X=341620 $Y=1101820
X79 694 1 2 18 BUF1S $T=350920 1112280 1 0 $X=350920 $Y=1106860
X80 30 1 2 56 BUF1S $T=419740 1092120 1 0 $X=419740 $Y=1086700
X81 56 1 2 48 BUF1S $T=422220 1102200 0 180 $X=419740 $Y=1096780
X82 59 1 2 55 BUF1S $T=429040 1122360 1 180 $X=426560 $Y=1121980
X83 57 1 2 765 BUF1S $T=442680 1102200 0 0 $X=442680 $Y=1101820
X84 129 1 2 144 BUF1S $T=501580 1092120 1 0 $X=501580 $Y=1086700
X85 144 1 2 169 BUF1S $T=526380 1112280 1 0 $X=526380 $Y=1106860
X86 170 1 2 166 BUF1S $T=531960 1112280 0 180 $X=529480 $Y=1106860
X87 166 1 2 196 BUF1S $T=553040 1092120 0 0 $X=553040 $Y=1091740
X88 841 1 2 205 BUF1S $T=579080 1112280 1 0 $X=579080 $Y=1106860
X89 205 1 2 223 BUF1S $T=590240 1092120 1 0 $X=590240 $Y=1086700
X90 869 1 2 886 BUF1S $T=604500 1112280 0 0 $X=604500 $Y=1111900
X91 248 1 2 896 BUF1S $T=617520 1102200 1 180 $X=615040 $Y=1101820
X92 250 1 2 244 BUF1S $T=619380 1092120 1 180 $X=616900 $Y=1091740
X93 886 1 2 915 BUF1S $T=636120 1122360 1 0 $X=636120 $Y=1116940
X94 266 1 2 881 BUF1S $T=647900 1102200 0 180 $X=645420 $Y=1096780
X95 276 1 2 893 BUF1S $T=657820 1092120 0 0 $X=657820 $Y=1091740
X96 299 1 2 968 BUF1S $T=691920 1102200 0 180 $X=689440 $Y=1096780
X97 299 1 2 983 BUF1S $T=703700 1092120 0 0 $X=703700 $Y=1091740
X98 968 1 2 989 BUF1S $T=708040 1122360 1 0 $X=708040 $Y=1116940
X99 316 1 2 283 BUF1S $T=734700 1092120 0 180 $X=732220 $Y=1086700
X100 319 1 2 315 BUF1S $T=740280 1092120 0 180 $X=737800 $Y=1086700
X101 982 1 2 1029 BUF1S $T=750200 1112280 0 0 $X=750200 $Y=1111900
X102 1026 1 2 1037 BUF1S $T=756400 1102200 1 0 $X=756400 $Y=1096780
X103 1035 1 2 1030 BUF1S $T=756400 1122360 1 0 $X=756400 $Y=1116940
X104 334 1 2 320 BUF1S $T=768800 1092120 1 180 $X=766320 $Y=1091740
X105 1098 1 2 1101 BUF1S $T=828940 1102200 0 0 $X=828940 $Y=1101820
X106 376 1 2 1099 BUF1S $T=839480 1102200 0 180 $X=837000 $Y=1096780
X107 1039 1 2 377 BUF1S $T=837620 1092120 0 0 $X=837620 $Y=1091740
X108 386 1 2 1127 BUF1S $T=852500 1102200 0 0 $X=852500 $Y=1101820
X109 1142 1 2 1144 BUF1S $T=867380 1122360 0 0 $X=867380 $Y=1121980
X110 1159 1 2 1176 BUF1S $T=896520 1112280 0 0 $X=896520 $Y=1111900
X111 1165 1 2 1182 BUF1S $T=908300 1102200 1 0 $X=908300 $Y=1096780
X112 1186 1 2 1193 BUF1S $T=928760 1102200 0 0 $X=928760 $Y=1101820
X113 447 1 2 438 BUF1S $T=934340 1092120 1 0 $X=934340 $Y=1086700
X114 452 1 2 450 BUF1S $T=943020 1092120 0 180 $X=940540 $Y=1086700
X115 452 1 2 1211 BUF1S $T=943640 1102200 0 0 $X=943640 $Y=1101820
X116 1208 1 2 1216 BUF1S $T=946740 1112280 0 0 $X=946740 $Y=1111900
X117 417 1 2 1197 BUF1S $T=961620 1112280 0 0 $X=961620 $Y=1111900
X118 1221 1 2 1229 BUF1S $T=964720 1102200 0 0 $X=964720 $Y=1101820
X119 493 1 2 1239 BUF1S $T=986420 1102200 1 0 $X=986420 $Y=1096780
X120 500 1 2 1204 BUF1S $T=993240 1102200 1 0 $X=993240 $Y=1096780
X121 428 1 2 521 BUF1S $T=1011220 1112280 0 0 $X=1011220 $Y=1111900
X122 475 1 2 520 BUF1S $T=1011840 1092120 1 0 $X=1011840 $Y=1086700
X123 524 1 2 1260 BUF1S $T=1023000 1102200 1 0 $X=1023000 $Y=1096780
X124 1260 1 2 1286 BUF1S $T=1037880 1122360 1 0 $X=1037880 $Y=1116940
X125 1338 1 2 651 BUF1S $T=1126540 1122360 0 0 $X=1126540 $Y=1121980
X126 682 1 2 683 DELB $T=291400 1092120 1 0 $X=291400 $Y=1086700
X127 687 1 2 688 DELB $T=308140 1112280 1 0 $X=308140 $Y=1106860
X128 696 1 2 15 DELB $T=329840 1092120 0 0 $X=329840 $Y=1091740
X129 699 1 2 700 DELB $T=332320 1112280 1 0 $X=332320 $Y=1106860
X130 702 1 2 705 DELB $T=336660 1102200 0 0 $X=336660 $Y=1101820
X131 23 1 2 28 DELB $T=345960 1102200 1 0 $X=345960 $Y=1096780
X132 715 1 2 718 DELB $T=355260 1102200 0 0 $X=355260 $Y=1101820
X133 716 1 2 717 DELB $T=362080 1092120 0 0 $X=362080 $Y=1091740
X134 727 1 2 733 DELB $T=393700 1122360 1 0 $X=393700 $Y=1116940
X135 729 1 2 738 DELB $T=399900 1112280 1 0 $X=399900 $Y=1106860
X136 739 1 2 742 DELB $T=406100 1112280 1 0 $X=406100 $Y=1106860
X137 746 1 2 748 DELB $T=412920 1112280 1 0 $X=412920 $Y=1106860
X138 752 1 2 751 DELB $T=422220 1092120 1 0 $X=422220 $Y=1086700
X139 756 1 2 758 DELB $T=426560 1102200 1 0 $X=426560 $Y=1096780
X140 67 1 2 71 DELB $T=435860 1092120 1 0 $X=435860 $Y=1086700
X141 760 1 2 764 DELB $T=443300 1092120 1 0 $X=443300 $Y=1086700
X142 82 1 2 86 DELB $T=450740 1092120 1 0 $X=450740 $Y=1086700
X143 774 1 2 773 DELB $T=454460 1112280 0 0 $X=454460 $Y=1111900
X144 92 1 2 95 DELB $T=461280 1112280 0 0 $X=461280 $Y=1111900
X145 785 1 2 786 DELB $T=466860 1092120 0 0 $X=466860 $Y=1091740
X146 791 1 2 793 DELB $T=471820 1112280 0 0 $X=471820 $Y=1111900
X147 107 1 2 116 DELB $T=475540 1102200 1 0 $X=475540 $Y=1096780
X148 801 1 2 799 DELB $T=488560 1112280 0 0 $X=488560 $Y=1111900
X149 804 1 2 803 DELB $T=491660 1092120 0 0 $X=491660 $Y=1091740
X150 807 1 2 808 DELB $T=496620 1112280 1 0 $X=496620 $Y=1106860
X151 809 1 2 810 DELB $T=497860 1092120 0 0 $X=497860 $Y=1091740
X152 813 1 2 818 DELB $T=505300 1092120 1 0 $X=505300 $Y=1086700
X153 816 1 2 817 DELB $T=507780 1112280 1 0 $X=507780 $Y=1106860
X154 152 1 2 158 DELB $T=512740 1092120 1 0 $X=512740 $Y=1086700
X155 820 1 2 819 DELB $T=512740 1112280 0 0 $X=512740 $Y=1111900
X156 156 1 2 162 DELB $T=515840 1122360 0 0 $X=515840 $Y=1121980
X157 823 1 2 827 DELB $T=517700 1092120 0 0 $X=517700 $Y=1091740
X158 831 1 2 832 DELB $T=532580 1122360 1 0 $X=532580 $Y=1116940
X159 835 1 2 834 DELB $T=538160 1092120 0 0 $X=538160 $Y=1091740
X160 185 1 2 191 DELB $T=544980 1102200 1 0 $X=544980 $Y=1096780
X161 844 1 2 845 DELB $T=553040 1102200 1 0 $X=553040 $Y=1096780
X162 199 1 2 202 DELB $T=556760 1122360 0 0 $X=556760 $Y=1121980
X163 848 1 2 843 DELB $T=558620 1092120 0 0 $X=558620 $Y=1091740
X164 855 1 2 852 DELB $T=565440 1122360 1 0 $X=565440 $Y=1116940
X165 851 1 2 857 DELB $T=566060 1092120 0 0 $X=566060 $Y=1091740
X166 211 1 2 216 DELB $T=571640 1122360 1 0 $X=571640 $Y=1116940
X167 859 1 2 860 DELB $T=572260 1102200 1 0 $X=572260 $Y=1096780
X168 854 1 2 862 DELB $T=574740 1112280 0 0 $X=574740 $Y=1111900
X169 861 1 2 864 DELB $T=579700 1092120 0 0 $X=579700 $Y=1091740
X170 221 1 2 224 DELB $T=581560 1112280 1 0 $X=581560 $Y=1106860
X171 222 1 2 873 DELB $T=585280 1092120 0 0 $X=585280 $Y=1091740
X172 889 1 2 891 DELB $T=610080 1112280 1 0 $X=610080 $Y=1106860
X173 895 1 2 894 DELB $T=611320 1122360 0 0 $X=611320 $Y=1121980
X174 903 1 2 907 DELB $T=618760 1122360 0 0 $X=618760 $Y=1121980
X175 901 1 2 911 DELB $T=624960 1102200 1 0 $X=624960 $Y=1096780
X176 902 1 2 912 DELB $T=633020 1102200 0 0 $X=633020 $Y=1101820
X177 919 1 2 923 DELB $T=642940 1122360 0 0 $X=642940 $Y=1121980
X178 270 1 2 274 DELB $T=651620 1122360 0 0 $X=651620 $Y=1121980
X179 935 1 2 936 DELB $T=652240 1102200 0 0 $X=652240 $Y=1101820
X180 937 1 2 934 DELB $T=653480 1122360 1 0 $X=653480 $Y=1116940
X181 941 1 2 933 DELB $T=660300 1092120 0 0 $X=660300 $Y=1091740
X182 940 1 2 946 DELB $T=660920 1122360 1 0 $X=660920 $Y=1116940
X183 280 1 2 282 DELB $T=666500 1092120 0 0 $X=666500 $Y=1091740
X184 950 1 2 954 DELB $T=669600 1122360 1 0 $X=669600 $Y=1116940
X185 286 1 2 290 DELB $T=677040 1122360 1 0 $X=677040 $Y=1116940
X186 287 1 2 292 DELB $T=678280 1092120 0 0 $X=678280 $Y=1091740
X187 958 1 2 957 DELB $T=681380 1112280 0 0 $X=681380 $Y=1111900
X188 965 1 2 970 DELB $T=690060 1112280 0 0 $X=690060 $Y=1111900
X189 972 1 2 975 DELB $T=695020 1122360 1 0 $X=695020 $Y=1116940
X190 991 1 2 998 DELB $T=716720 1102200 1 0 $X=716720 $Y=1096780
X191 1001 1 2 1010 DELB $T=722920 1102200 1 0 $X=722920 $Y=1096780
X192 1003 1 2 1006 DELB $T=726020 1122360 1 0 $X=726020 $Y=1116940
X193 1009 1 2 1015 DELB $T=727260 1092120 1 0 $X=727260 $Y=1086700
X194 324 1 2 327 DELB $T=750820 1102200 1 0 $X=750820 $Y=1096780
X195 330 1 2 332 DELB $T=758880 1102200 1 0 $X=758880 $Y=1096780
X196 336 1 2 340 DELB $T=776860 1092120 1 0 $X=776860 $Y=1086700
X197 339 1 2 342 DELB $T=778100 1122360 0 0 $X=778100 $Y=1121980
X198 1063 1 2 1066 DELB $T=782440 1102200 0 0 $X=782440 $Y=1101820
X199 1067 1 2 1068 DELB $T=786160 1122360 0 0 $X=786160 $Y=1121980
X200 349 1 2 353 DELB $T=791120 1092120 1 0 $X=791120 $Y=1086700
X201 1075 1 2 1079 DELB $T=794220 1122360 0 0 $X=794220 $Y=1121980
X202 1074 1 2 1065 DELB $T=795460 1102200 1 0 $X=795460 $Y=1096780
X203 355 1 2 358 DELB $T=800420 1112280 1 0 $X=800420 $Y=1106860
X204 1087 1 2 1085 DELB $T=804140 1092120 0 0 $X=804140 $Y=1091740
X205 364 1 2 367 DELB $T=814680 1122360 0 0 $X=814680 $Y=1121980
X206 368 1 2 370 DELB $T=821500 1122360 0 0 $X=821500 $Y=1121980
X207 1094 1 2 1104 DELB $T=822740 1112280 1 0 $X=822740 $Y=1106860
X208 1096 1 2 1105 DELB $T=827700 1112280 0 0 $X=827700 $Y=1111900
X209 1118 1 2 1124 DELB $T=844440 1112280 1 0 $X=844440 $Y=1106860
X210 1129 1 2 1137 DELB $T=852500 1112280 0 0 $X=852500 $Y=1111900
X211 1148 1 2 1152 DELB $T=869240 1112280 0 0 $X=869240 $Y=1111900
X212 1145 1 2 1154 DELB $T=875440 1112280 1 0 $X=875440 $Y=1106860
X213 1161 1 2 1167 DELB $T=887220 1102200 1 0 $X=887220 $Y=1096780
X214 421 1 2 425 DELB $T=903960 1102200 0 0 $X=903960 $Y=1101820
X215 1044 1 2 1043 DELB $T=917600 1122360 0 0 $X=917600 $Y=1121980
X216 431 1 2 440 DELB $T=920700 1112280 0 0 $X=920700 $Y=1111900
X217 446 1 2 449 DELB $T=934340 1122360 0 0 $X=934340 $Y=1121980
X218 1219 1 2 1224 DELB $T=955420 1112280 1 0 $X=955420 $Y=1106860
X219 467 1 2 472 DELB $T=958520 1092120 1 0 $X=958520 $Y=1086700
X220 1222 1 2 1223 DELB $T=959140 1102200 0 0 $X=959140 $Y=1101820
X221 470 1 2 477 DELB $T=959760 1122360 0 0 $X=959760 $Y=1121980
X222 1228 1 2 1231 DELB $T=967820 1102200 0 0 $X=967820 $Y=1101820
X223 487 1 2 490 DELB $T=974640 1112280 0 0 $X=974640 $Y=1111900
X224 492 1 2 496 DELB $T=983320 1112280 0 0 $X=983320 $Y=1111900
X225 1254 1 2 1253 DELB $T=1001300 1092120 0 0 $X=1001300 $Y=1091740
X226 1262 1 2 1267 DELB $T=1008120 1092120 0 0 $X=1008120 $Y=1091740
X227 1269 1 2 1273 DELB $T=1018040 1112280 0 0 $X=1018040 $Y=1111900
X228 1277 1 2 1276 DELB $T=1027960 1112280 0 0 $X=1027960 $Y=1111900
X229 544 1 2 550 DELB $T=1040360 1122360 1 0 $X=1040360 $Y=1116940
X230 1279 1 2 1282 DELB $T=1042840 1112280 1 0 $X=1042840 $Y=1106860
X231 590 1 2 595 DELB $T=1080040 1092120 1 0 $X=1080040 $Y=1086700
X232 546 1 2 1295 DELB $T=1080660 1112280 1 0 $X=1080660 $Y=1106860
X233 598 1 2 603 DELB $T=1085000 1122360 0 0 $X=1085000 $Y=1121980
X234 1316 1 2 1317 DELB $T=1086860 1092120 1 0 $X=1086860 $Y=1086700
X235 1318 1 2 1319 DELB $T=1089960 1102200 0 0 $X=1089960 $Y=1101820
X236 1328 1 2 1327 DELB $T=1099880 1112280 1 0 $X=1099880 $Y=1106860
X237 619 1 2 625 DELB $T=1105460 1102200 1 0 $X=1105460 $Y=1096780
X238 1332 1 2 1333 DELB $T=1110420 1092120 0 0 $X=1110420 $Y=1091740
X239 643 1 2 648 DELB $T=1121580 1122360 0 0 $X=1121580 $Y=1121980
X240 644 1 2 650 DELB $T=1122200 1112280 0 0 $X=1122200 $Y=1111900
X241 63 1 2 68 DELA $T=431520 1122360 1 0 $X=431520 $Y=1116940
X242 72 1 2 78 DELA $T=441440 1122360 0 0 $X=441440 $Y=1121980
X243 99 1 2 103 DELA $T=466240 1122360 0 0 $X=466240 $Y=1121980
X244 100 1 2 104 DELA $T=466860 1112280 0 0 $X=466860 $Y=1111900
X245 119 1 2 124 DELA $T=481120 1122360 0 0 $X=481120 $Y=1121980
X246 123 1 2 131 DELA $T=484220 1122360 1 0 $X=484220 $Y=1116940
X247 163 1 2 167 DELA $T=522040 1122360 0 0 $X=522040 $Y=1121980
X248 168 1 2 172 DELA $T=527000 1122360 0 0 $X=527000 $Y=1121980
X249 195 1 2 198 DELA $T=551800 1122360 0 0 $X=551800 $Y=1121980
X250 215 1 2 218 DELA $T=572880 1122360 0 0 $X=572880 $Y=1121980
X251 227 1 2 230 DELA $T=591480 1122360 0 0 $X=591480 $Y=1121980
X252 231 1 2 235 DELA $T=596440 1122360 0 0 $X=596440 $Y=1121980
X253 253 1 2 254 DELA $T=628060 1122360 0 0 $X=628060 $Y=1121980
X254 255 1 2 260 DELA $T=633020 1122360 0 0 $X=633020 $Y=1121980
X255 261 1 2 265 DELA $T=637980 1122360 0 0 $X=637980 $Y=1121980
X256 344 1 2 347 DELA $T=786160 1092120 1 0 $X=786160 $Y=1086700
X257 427 1 2 430 DELA $T=912640 1122360 0 0 $X=912640 $Y=1121980
X258 457 1 2 462 DELA $T=948600 1092120 1 0 $X=948600 $Y=1086700
X259 460 1 2 466 DELA $T=951700 1122360 0 0 $X=951700 $Y=1121980
X260 497 1 2 502 DELA $T=987660 1122360 1 0 $X=987660 $Y=1116940
X261 507 1 2 512 DELA $T=999440 1122360 0 0 $X=999440 $Y=1121980
X262 533 1 2 537 DELA $T=1030440 1122360 0 0 $X=1030440 $Y=1121980
X263 539 1 2 545 DELA $T=1036640 1122360 0 0 $X=1036640 $Y=1121980
X264 548 1 2 556 DELA $T=1045320 1122360 0 0 $X=1045320 $Y=1121980
X265 566 1 2 572 DELA $T=1060200 1122360 0 0 $X=1060200 $Y=1121980
X266 596 1 2 602 DELA $T=1084380 1102200 0 0 $X=1084380 $Y=1101820
X267 613 1 2 618 DELA $T=1100500 1102200 1 0 $X=1100500 $Y=1096780
X268 614 1 2 620 DELA $T=1101120 1122360 1 0 $X=1101120 $Y=1116940
X269 616 1 2 622 DELA $T=1101740 1122360 0 0 $X=1101740 $Y=1121980
X270 621 1 2 626 DELA $T=1106080 1122360 1 0 $X=1106080 $Y=1116940
X271 628 1 2 631 DELA $T=1111040 1122360 1 0 $X=1111040 $Y=1116940
X272 632 1 2 638 DELA $T=1116000 1122360 1 0 $X=1116000 $Y=1116940
X273 635 1 2 641 DELA $T=1116620 1122360 0 0 $X=1116620 $Y=1121980
X274 640 1 2 646 DELA $T=1120960 1122360 1 0 $X=1120960 $Y=1116940
X275 642 1 2 647 DELA $T=1121580 1112280 1 0 $X=1121580 $Y=1106860
X276 683 7 5 2 1 686 QDFFRBN $T=292640 1092120 0 0 $X=292640 $Y=1091740
X277 688 7 694 2 1 690 QDFFRBN $T=307520 1102200 0 0 $X=307520 $Y=1101820
X278 11 7 5 2 1 14 QDFFRBN $T=308140 1092120 1 0 $X=308140 $Y=1086700
X279 700 7 694 2 1 689 QDFFRBN $T=334180 1102200 1 180 $X=322400 $Y=1101820
X280 16 7 18 2 1 696 QDFFRBN $T=326120 1092120 1 0 $X=326120 $Y=1086700
X281 703 7 18 2 1 702 QDFFRBN $T=337280 1112280 1 0 $X=337280 $Y=1106860
X282 717 7 18 2 1 21 QDFFRBN $T=367040 1092120 0 180 $X=355260 $Y=1086700
X283 718 7 694 2 1 714 QDFFRBN $T=368900 1102200 0 180 $X=357120 $Y=1096780
X284 719 32 722 2 1 725 QDFFRBN $T=370140 1102200 0 0 $X=370140 $Y=1101820
X285 720 32 722 2 1 33 QDFFRBN $T=371380 1092120 1 0 $X=371380 $Y=1086700
X286 721 32 722 2 1 726 QDFFRBN $T=372000 1102200 1 0 $X=372000 $Y=1096780
X287 723 32 722 2 1 727 QDFFRBN $T=373860 1112280 1 0 $X=373860 $Y=1106860
X288 736 32 722 2 1 729 QDFFRBN $T=401140 1112280 1 180 $X=389360 $Y=1111900
X289 734 32 48 2 1 47 QDFFRBN $T=394320 1092120 0 0 $X=394320 $Y=1091740
X290 740 32 48 2 1 739 QDFFRBN $T=402380 1102200 0 0 $X=402380 $Y=1101820
X291 741 32 48 2 1 746 QDFFRBN $T=404240 1112280 0 0 $X=404240 $Y=1111900
X292 743 32 48 2 1 752 QDFFRBN $T=407340 1092120 0 0 $X=407340 $Y=1091740
X293 750 32 48 2 1 756 QDFFRBN $T=417880 1112280 1 0 $X=417880 $Y=1106860
X294 761 61 56 2 1 755 QDFFRBN $T=434000 1092120 1 180 $X=422220 $Y=1091740
X295 766 61 722 2 1 759 QDFFRBN $T=443920 1112280 0 180 $X=432140 $Y=1106860
X296 762 61 767 2 1 760 QDFFRBN $T=435860 1102200 1 0 $X=435860 $Y=1096780
X297 85 61 76 2 1 64 QDFFRBN $T=454460 1092120 1 180 $X=442680 $Y=1091740
X298 768 61 767 2 1 771 QDFFRBN $T=446400 1112280 1 0 $X=446400 $Y=1106860
X299 769 61 767 2 1 774 QDFFRBN $T=446400 1122360 1 0 $X=446400 $Y=1116940
X300 772 61 767 2 1 781 QDFFRBN $T=450120 1102200 1 0 $X=450120 $Y=1096780
X301 780 61 767 2 1 785 QDFFRBN $T=461280 1112280 1 0 $X=461280 $Y=1106860
X302 782 61 789 2 1 791 QDFFRBN $T=461900 1122360 1 0 $X=461900 $Y=1116940
X303 94 61 767 2 1 776 QDFFRBN $T=463760 1102200 1 0 $X=463760 $Y=1096780
X304 795 61 789 2 1 801 QDFFRBN $T=476780 1112280 0 0 $X=476780 $Y=1111900
X305 800 61 118 2 1 109 QDFFRBN $T=489800 1092120 1 180 $X=478020 $Y=1091740
X306 797 61 789 2 1 804 QDFFRBN $T=481120 1102200 0 0 $X=481120 $Y=1101820
X307 802 61 789 2 1 807 QDFFRBN $T=489180 1122360 1 0 $X=489180 $Y=1116940
X308 805 61 118 2 1 809 QDFFRBN $T=491660 1102200 1 0 $X=491660 $Y=1096780
X309 806 61 789 2 1 816 QDFFRBN $T=493520 1112280 0 0 $X=493520 $Y=1111900
X310 814 61 789 2 1 820 QDFFRBN $T=504060 1122360 1 0 $X=504060 $Y=1116940
X311 815 61 153 2 1 155 QDFFRBN $T=504680 1092120 0 0 $X=504680 $Y=1091740
X312 812 61 153 2 1 813 QDFFRBN $T=505300 1102200 1 0 $X=505300 $Y=1096780
X313 824 61 166 2 1 823 QDFFRBN $T=517080 1102200 0 0 $X=517080 $Y=1101820
X314 826 61 166 2 1 825 QDFFRBN $T=517700 1112280 0 0 $X=517700 $Y=1111900
X315 829 61 170 2 1 835 QDFFRBN $T=525760 1092120 1 0 $X=525760 $Y=1086700
X316 839 182 170 2 1 830 QDFFRBN $T=543120 1102200 1 180 $X=531340 $Y=1101820
X317 833 61 166 2 1 831 QDFFRBN $T=532580 1112280 0 0 $X=532580 $Y=1111900
X318 838 182 170 2 1 174 QDFFRBN $T=544980 1102200 0 180 $X=533200 $Y=1096780
X319 186 182 196 2 1 197 QDFFRBN $T=544980 1092120 1 0 $X=544980 $Y=1086700
X320 840 182 166 2 1 848 QDFFRBN $T=545600 1102200 0 0 $X=545600 $Y=1101820
X321 842 182 841 2 1 844 QDFFRBN $T=547460 1112280 0 0 $X=547460 $Y=1111900
X322 846 182 841 2 1 855 QDFFRBN $T=553660 1122360 1 0 $X=553660 $Y=1116940
X323 201 182 205 2 1 106 QDFFRBN $T=558620 1092120 1 0 $X=558620 $Y=1086700
X324 850 182 205 2 1 851 QDFFRBN $T=558620 1102200 0 0 $X=558620 $Y=1101820
X325 863 182 841 2 1 854 QDFFRBN $T=574740 1112280 1 180 $X=562960 $Y=1111900
X326 872 182 869 2 1 853 QDFFRBN $T=588380 1122360 0 180 $X=576600 $Y=1116940
X327 220 182 223 2 1 226 QDFFRBN $T=577840 1092120 1 0 $X=577840 $Y=1086700
X328 865 182 205 2 1 859 QDFFRBN $T=590240 1102200 1 180 $X=578460 $Y=1101820
X329 868 182 225 2 1 861 QDFFRBN $T=579700 1102200 1 0 $X=579700 $Y=1096780
X330 882 182 869 2 1 874 QDFFRBN $T=602020 1092120 1 180 $X=590240 $Y=1091740
X331 875 182 869 2 1 879 QDFFRBN $T=590240 1112280 0 0 $X=590240 $Y=1111900
X332 877 182 869 2 1 883 QDFFRBN $T=591480 1122360 1 0 $X=591480 $Y=1116940
X333 878 182 225 2 1 889 QDFFRBN $T=595200 1102200 1 0 $X=595200 $Y=1096780
X334 234 182 225 2 1 242 QDFFRBN $T=599540 1092120 1 0 $X=599540 $Y=1086700
X335 887 182 886 2 1 895 QDFFRBN $T=606360 1122360 1 0 $X=606360 $Y=1116940
X336 900 182 886 2 1 903 QDFFRBN $T=614420 1112280 0 0 $X=614420 $Y=1111900
X337 914 182 252 2 1 901 QDFFRBN $T=633020 1092120 0 180 $X=621240 $Y=1086700
X338 908 182 886 2 1 866 QDFFRBN $T=621240 1122360 1 0 $X=621240 $Y=1116940
X339 910 182 915 2 1 902 QDFFRBN $T=621860 1112280 1 0 $X=621860 $Y=1106860
X340 913 182 886 2 1 919 QDFFRBN $T=628680 1112280 0 0 $X=628680 $Y=1111900
X341 916 182 262 2 1 920 QDFFRBN $T=631160 1092120 0 0 $X=631160 $Y=1091740
X342 917 182 915 2 1 924 QDFFRBN $T=635500 1112280 1 0 $X=635500 $Y=1106860
X343 922 182 915 2 1 937 QDFFRBN $T=641700 1122360 1 0 $X=641700 $Y=1116940
X344 927 182 262 2 1 941 QDFFRBN $T=645420 1092120 0 0 $X=645420 $Y=1091740
X345 939 279 915 2 1 935 QDFFRBN $T=668360 1122360 1 180 $X=656580 $Y=1121980
X346 948 279 915 2 1 940 QDFFRBN $T=668980 1112280 1 180 $X=657200 $Y=1111900
X347 949 279 915 2 1 942 QDFFRBN $T=669600 1102200 1 180 $X=657820 $Y=1101820
X348 278 182 281 2 1 284 QDFFRBN $T=660300 1092120 1 0 $X=660300 $Y=1086700
X349 956 279 281 2 1 950 QDFFRBN $T=680760 1112280 0 180 $X=668980 $Y=1106860
X350 951 279 281 2 1 958 QDFFRBN $T=670840 1122360 0 0 $X=670840 $Y=1121980
X351 963 279 281 2 1 955 QDFFRBN $T=685720 1102200 1 180 $X=673940 $Y=1101820
X352 285 182 281 2 1 287 QDFFRBN $T=675180 1092120 1 0 $X=675180 $Y=1086700
X353 967 279 281 2 1 959 QDFFRBN $T=693780 1122360 0 180 $X=682000 $Y=1116940
X354 964 279 968 2 1 972 QDFFRBN $T=685720 1122360 0 0 $X=685720 $Y=1121980
X355 973 279 968 2 1 965 QDFFRBN $T=699360 1102200 1 180 $X=687580 $Y=1101820
X356 297 182 299 2 1 304 QDFFRBN $T=690060 1092120 0 0 $X=690060 $Y=1091740
X357 302 182 983 2 1 305 QDFFRBN $T=699360 1092120 1 0 $X=699360 $Y=1086700
X358 978 279 968 2 1 985 QDFFRBN $T=700600 1122360 0 0 $X=700600 $Y=1121980
X359 979 279 983 2 1 306 QDFFRBN $T=701220 1102200 1 0 $X=701220 $Y=1096780
X360 984 279 968 2 1 980 QDFFRBN $T=713620 1102200 1 180 $X=701840 $Y=1101820
X361 310 279 983 2 1 307 QDFFRBN $T=725400 1092120 0 180 $X=713620 $Y=1086700
X362 1005 279 983 2 1 993 QDFFRBN $T=726020 1092120 1 180 $X=714240 $Y=1091740
X363 999 279 983 2 1 991 QDFFRBN $T=726640 1102200 1 180 $X=714860 $Y=1101820
X364 1000 279 989 2 1 996 QDFFRBN $T=727260 1122360 1 180 $X=715480 $Y=1121980
X365 1020 279 989 2 1 1011 QDFFRBN $T=739660 1102200 1 180 $X=727880 $Y=1101820
X366 1013 279 989 2 1 1003 QDFFRBN $T=741520 1122360 1 180 $X=729740 $Y=1121980
X367 1022 279 989 2 1 1014 QDFFRBN $T=744620 1122360 0 180 $X=732840 $Y=1116940
X368 1019 279 989 2 1 1001 QDFFRBN $T=750820 1102200 0 180 $X=739040 $Y=1096780
X369 1027 279 320 2 1 1009 QDFFRBN $T=752680 1092120 1 180 $X=740900 $Y=1091740
X370 1025 279 989 2 1 1007 QDFFRBN $T=753920 1102200 1 180 $X=742140 $Y=1101820
X371 1024 279 320 2 1 1035 QDFFRBN $T=744620 1122360 0 0 $X=744620 $Y=1121980
X372 1031 279 320 2 1 1026 QDFFRBN $T=761360 1092120 0 180 $X=749580 $Y=1086700
X373 1033 279 320 2 1 1044 QDFFRBN $T=755160 1102200 0 0 $X=755160 $Y=1101820
X374 1034 279 320 2 1 1040 QDFFRBN $T=755160 1112280 1 0 $X=755160 $Y=1106860
X375 1038 279 1045 2 1 1046 QDFFRBN $T=758880 1122360 1 0 $X=758880 $Y=1116940
X376 1051 279 334 2 1 1042 QDFFRBN $T=776860 1092120 0 180 $X=765080 $Y=1086700
X377 1049 279 1045 2 1 1052 QDFFRBN $T=768800 1112280 1 0 $X=768800 $Y=1106860
X378 1050 341 1045 2 1 1053 QDFFRBN $T=784920 1122360 0 180 $X=773140 $Y=1116940
X379 1059 279 334 2 1 1074 QDFFRBN $T=778720 1092120 0 0 $X=778720 $Y=1091740
X380 1062 279 1073 2 1 1063 QDFFRBN $T=783060 1112280 1 0 $X=783060 $Y=1106860
X381 1064 341 1073 2 1 1067 QDFFRBN $T=786780 1122360 1 0 $X=786780 $Y=1116940
X382 1080 341 351 2 1 1075 QDFFRBN $T=803520 1102200 1 180 $X=791740 $Y=1101820
X383 1082 341 351 2 1 1087 QDFFRBN $T=799180 1092120 1 0 $X=799180 $Y=1086700
X384 1083 341 1073 2 1 1093 QDFFRBN $T=800420 1122360 1 0 $X=800420 $Y=1116940
X385 1084 341 1073 2 1 1091 QDFFRBN $T=802900 1122360 0 0 $X=802900 $Y=1121980
X386 1086 341 1073 2 1 360 QDFFRBN $T=803520 1102200 0 0 $X=803520 $Y=1101820
X387 1100 341 351 2 1 361 QDFFRBN $T=824600 1092120 0 180 $X=812820 $Y=1086700
X388 1106 341 351 2 1 1089 QDFFRBN $T=825840 1102200 0 180 $X=814060 $Y=1096780
X389 1095 341 1099 2 1 1094 QDFFRBN $T=815300 1122360 1 0 $X=815300 $Y=1116940
X390 1107 341 1099 2 1 1096 QDFFRBN $T=828940 1102200 1 180 $X=817160 $Y=1101820
X391 1113 341 1099 2 1 1098 QDFFRBN $T=838240 1122360 1 180 $X=826460 $Y=1121980
X392 1108 341 372 2 1 375 QDFFRBN $T=827080 1092120 1 0 $X=827080 $Y=1086700
X393 1111 341 1099 2 1 1117 QDFFRBN $T=830800 1122360 1 0 $X=830800 $Y=1116940
X394 1120 341 1099 2 1 1112 QDFFRBN $T=843200 1102200 1 180 $X=831420 $Y=1101820
X395 378 341 376 2 1 379 QDFFRBN $T=840100 1092120 0 0 $X=840100 $Y=1091740
X396 1121 341 376 2 1 1118 QDFFRBN $T=852500 1102200 0 180 $X=840720 $Y=1096780
X397 1119 341 1099 2 1 1122 QDFFRBN $T=840720 1122360 0 0 $X=840720 $Y=1121980
X398 388 341 1142 2 1 394 QDFFRBN $T=853120 1092120 1 0 $X=853120 $Y=1086700
X399 1133 341 1142 2 1 1143 QDFFRBN $T=854360 1102200 1 0 $X=854360 $Y=1096780
X400 1134 341 1142 2 1 1132 QDFFRBN $T=854360 1122360 1 0 $X=854360 $Y=1116940
X401 1139 341 1144 2 1 1129 QDFFRBN $T=857460 1112280 0 0 $X=857460 $Y=1111900
X402 1155 341 1142 2 1 400 QDFFRBN $T=880400 1092120 1 180 $X=868620 $Y=1091740
X403 1157 341 1142 2 1 1145 QDFFRBN $T=880400 1102200 0 180 $X=868620 $Y=1096780
X404 1149 341 1144 2 1 1148 QDFFRBN $T=869860 1122360 1 0 $X=869860 $Y=1116940
X405 1170 411 1165 2 1 1161 QDFFRBN $T=894660 1092120 1 180 $X=882880 $Y=1091740
X406 1158 341 1144 2 1 1160 QDFFRBN $T=895280 1122360 0 180 $X=883500 $Y=1116940
X407 1163 341 1144 2 1 1169 QDFFRBN $T=884740 1112280 0 0 $X=884740 $Y=1111900
X408 1156 411 1165 2 1 1123 QDFFRBN $T=901480 1092120 0 180 $X=889700 $Y=1086700
X409 1178 411 1165 2 1 1166 QDFFRBN $T=905820 1102200 0 180 $X=894040 $Y=1096780
X410 1172 411 1144 2 1 1159 QDFFRBN $T=908920 1122360 0 180 $X=897140 $Y=1116940
X411 1180 411 1144 2 1 1171 QDFFRBN $T=910780 1112280 1 180 $X=899000 $Y=1111900
X412 1177 411 1165 2 1 1164 QDFFRBN $T=912640 1092120 1 180 $X=900860 $Y=1091740
X413 429 411 422 2 1 420 QDFFRBN $T=915740 1092120 0 180 $X=903960 $Y=1086700
X414 1181 411 1182 2 1 1188 QDFFRBN $T=908920 1102200 0 0 $X=908920 $Y=1101820
X415 1183 411 1182 2 1 1187 QDFFRBN $T=911400 1122360 1 0 $X=911400 $Y=1116940
X416 1184 411 1182 2 1 432 QDFFRBN $T=913260 1102200 1 0 $X=913260 $Y=1096780
X417 1191 411 1182 2 1 1186 QDFFRBN $T=930000 1112280 0 180 $X=918220 $Y=1106860
X418 1196 411 1182 2 1 439 QDFFRBN $T=933720 1092120 1 180 $X=921940 $Y=1091740
X419 1200 411 1182 2 1 1190 QDFFRBN $T=936200 1122360 0 180 $X=924420 $Y=1116940
X420 1202 411 1211 2 1 1205 QDFFRBN $T=934960 1112280 0 0 $X=934960 $Y=1111900
X421 1207 411 450 2 1 1199 QDFFRBN $T=947980 1092120 1 180 $X=936200 $Y=1091740
X422 1203 411 1211 2 1 1212 QDFFRBN $T=937440 1122360 1 0 $X=937440 $Y=1116940
X423 1220 411 452 2 1 1209 QDFFRBN $T=953560 1102200 0 180 $X=941780 $Y=1096780
X424 1215 411 1211 2 1 1222 QDFFRBN $T=946740 1102200 0 0 $X=946740 $Y=1101820
X425 1217 411 1211 2 1 1219 QDFFRBN $T=952320 1122360 1 0 $X=952320 $Y=1116940
X426 1225 411 1211 2 1 1228 QDFFRBN $T=960380 1112280 1 0 $X=960380 $Y=1106860
X427 486 411 452 2 1 473 QDFFRBN $T=975260 1092120 0 180 $X=963480 $Y=1086700
X428 1232 411 1211 2 1 1221 QDFFRBN $T=977120 1122360 1 180 $X=965340 $Y=1121980
X429 1235 411 1239 2 1 482 QDFFRBN $T=973400 1102200 1 0 $X=973400 $Y=1096780
X430 1234 411 1239 2 1 478 QDFFRBN $T=973400 1102200 0 0 $X=973400 $Y=1101820
X431 1237 411 1239 2 1 1240 QDFFRBN $T=974640 1112280 1 0 $X=974640 $Y=1106860
X432 1236 411 1239 2 1 1230 QDFFRBN $T=975880 1122360 1 0 $X=975880 $Y=1116940
X433 1238 411 493 2 1 498 QDFFRBN $T=977120 1092120 0 0 $X=977120 $Y=1091740
X434 489 411 493 2 1 499 QDFFRBN $T=977740 1092120 1 0 $X=977740 $Y=1086700
X435 1241 411 1239 2 1 1243 QDFFRBN $T=987040 1102200 0 0 $X=987040 $Y=1101820
X436 1242 411 1239 2 1 1249 QDFFRBN $T=987660 1122360 0 0 $X=987660 $Y=1121980
X437 1250 411 1260 2 1 1264 QDFFRBN $T=997580 1112280 0 0 $X=997580 $Y=1111900
X438 1247 411 493 2 1 1254 QDFFRBN $T=1011220 1102200 1 180 $X=999440 $Y=1101820
X439 1266 411 1260 2 1 1269 QDFFRBN $T=1008740 1122360 1 0 $X=1008740 $Y=1116940
X440 1271 527 524 2 1 1262 QDFFRBN $T=1024860 1092120 1 180 $X=1013080 $Y=1091740
X441 1270 411 524 2 1 1265 QDFFRBN $T=1014320 1112280 1 0 $X=1014320 $Y=1106860
X442 1268 527 1260 2 1 523 QDFFRBN $T=1027340 1092120 0 180 $X=1015560 $Y=1086700
X443 1274 527 1260 2 1 1277 QDFFRBN $T=1023620 1122360 1 0 $X=1023620 $Y=1116940
X444 1275 527 1260 2 1 1283 QDFFRBN $T=1027340 1102200 1 0 $X=1027340 $Y=1096780
X445 1281 527 1286 2 1 1285 QDFFRBN $T=1031680 1102200 0 0 $X=1031680 $Y=1101820
X446 1278 527 1286 2 1 1279 QDFFRBN $T=1033540 1112280 0 0 $X=1033540 $Y=1111900
X447 1293 527 555 2 1 549 QDFFRBN $T=1056480 1092120 1 180 $X=1044700 $Y=1091740
X448 1289 527 1286 2 1 1297 QDFFRBN $T=1045320 1102200 0 0 $X=1045320 $Y=1101820
X449 1288 527 1286 2 1 1291 QDFFRBN $T=1045320 1122360 1 0 $X=1045320 $Y=1116940
X450 1304 527 1286 2 1 1300 QDFFRBN $T=1070740 1102200 1 180 $X=1058960 $Y=1101820
X451 1302 527 569 2 1 552 QDFFRBN $T=1071360 1092120 1 180 $X=1059580 $Y=1091740
X452 1303 527 1286 2 1 1296 QDFFRBN $T=1075080 1112280 1 180 $X=1063300 $Y=1111900
X453 578 527 583 2 1 588 QDFFRBN $T=1068260 1092120 1 0 $X=1068260 $Y=1086700
X454 1312 527 583 2 1 1307 QDFFRBN $T=1082520 1102200 0 180 $X=1070740 $Y=1096780
X455 1315 527 1311 2 1 1308 QDFFRBN $T=1084380 1102200 1 180 $X=1072600 $Y=1101820
X456 1313 527 1311 2 1 1318 QDFFRBN $T=1078800 1112280 0 0 $X=1078800 $Y=1111900
X457 1314 527 1311 2 1 1316 QDFFRBN $T=1084380 1102200 1 0 $X=1084380 $Y=1096780
X458 1323 527 1311 2 1 1328 QDFFRBN $T=1094300 1112280 0 0 $X=1094300 $Y=1111900
X459 1320 527 583 2 1 601 QDFFRBN $T=1109800 1092120 0 180 $X=1098020 $Y=1086700
X460 1321 527 583 2 1 1326 QDFFRBN $T=1110420 1102200 1 180 $X=1098640 $Y=1101820
X461 1335 527 1311 2 1 1329 QDFFRBN $T=1122200 1112280 1 180 $X=1110420 $Y=1111900
X462 1336 527 1311 2 1 1330 QDFFRBN $T=1125920 1102200 1 180 $X=1114140 $Y=1101820
X463 649 527 636 2 1 624 QDFFRBN $T=1128400 1092120 0 180 $X=1116620 $Y=1086700
X464 1337 527 636 2 1 1332 QDFFRBN $T=1128400 1092120 1 180 $X=1116620 $Y=1091740
X465 33 1 2 724 34 35 681 ICV_4 $T=375720 1092120 0 0 $X=375720 $Y=1091740
X466 726 1 2 730 725 728 681 ICV_4 $T=389980 1112280 1 0 $X=389980 $Y=1106860
X467 64 1 2 69 759 763 681 ICV_4 $T=432140 1112280 0 0 $X=432140 $Y=1111900
X468 75 1 2 80 771 770 681 ICV_4 $T=444540 1112280 0 0 $X=444540 $Y=1111900
X469 79 1 2 83 84 87 681 ICV_4 $T=446400 1122360 0 0 $X=446400 $Y=1121980
X470 89 1 2 90 93 96 681 ICV_4 $T=456320 1122360 0 0 $X=456320 $Y=1121980
X471 776 1 2 91 781 783 681 ICV_4 $T=456940 1092120 0 0 $X=456940 $Y=1091740
X472 126 1 2 133 136 139 681 ICV_4 $T=486080 1122360 0 0 $X=486080 $Y=1121980
X473 140 1 2 142 143 145 681 ICV_4 $T=496000 1122360 0 0 $X=496000 $Y=1121980
X474 160 1 2 165 825 828 681 ICV_4 $T=520180 1122360 1 0 $X=520180 $Y=1116940
X475 830 1 2 837 187 192 681 ICV_4 $T=541260 1122360 1 0 $X=541260 $Y=1116940
X476 184 1 2 188 190 194 681 ICV_4 $T=541880 1122360 0 0 $X=541880 $Y=1121980
X477 203 1 2 208 209 212 681 ICV_4 $T=562960 1122360 0 0 $X=562960 $Y=1121980
X478 866 1 2 870 853 871 681 ICV_4 $T=577840 1122360 0 0 $X=577840 $Y=1121980
X479 879 1 2 880 883 884 681 ICV_4 $T=596440 1102200 0 0 $X=596440 $Y=1101820
X480 236 1 2 238 239 241 681 ICV_4 $T=601400 1122360 0 0 $X=601400 $Y=1121980
X481 242 1 2 247 874 890 681 ICV_4 $T=611320 1092120 1 0 $X=611320 $Y=1086700
X482 920 1 2 918 924 921 681 ICV_4 $T=641700 1102200 0 0 $X=641700 $Y=1101820
X483 942 1 2 947 284 288 681 ICV_4 $T=670840 1102200 1 0 $X=670840 $Y=1096780
X484 955 1 2 966 959 969 681 ICV_4 $T=688200 1092120 1 0 $X=688200 $Y=1086700
X485 980 1 2 981 985 986 681 ICV_4 $T=702460 1112280 0 0 $X=702460 $Y=1111900
X486 996 1 2 997 306 990 681 ICV_4 $T=716100 1122360 1 0 $X=716100 $Y=1116940
X487 993 1 2 1017 1011 1018 681 ICV_4 $T=729120 1112280 0 0 $X=729120 $Y=1111900
X488 1014 1 2 1021 322 325 681 ICV_4 $T=742760 1112280 1 0 $X=742760 $Y=1106860
X489 1007 1 2 1023 323 326 681 ICV_4 $T=744620 1122360 1 0 $X=744620 $Y=1116940
X490 328 1 2 331 1040 1041 681 ICV_4 $T=757640 1122360 0 0 $X=757640 $Y=1121980
X491 1042 1 2 1048 1052 1054 681 ICV_4 $T=768180 1102200 1 0 $X=768180 $Y=1096780
X492 1046 1 2 1047 1053 1055 681 ICV_4 $T=768180 1122360 0 0 $X=768180 $Y=1121980
X493 361 1 2 1097 1089 1102 681 ICV_4 $T=825840 1092120 0 0 $X=825840 $Y=1091740
X494 1112 1 2 1115 1117 1116 681 ICV_4 $T=834520 1112280 0 0 $X=834520 $Y=1111900
X495 379 1 2 382 1123 1128 681 ICV_4 $T=843200 1092120 1 0 $X=843200 $Y=1086700
X496 380 1 2 384 1122 1125 681 ICV_4 $T=843200 1122360 1 0 $X=843200 $Y=1116940
X497 1132 1 2 1131 1093 1088 681 ICV_4 $T=853120 1122360 0 0 $X=853120 $Y=1121980
X498 387 1 2 390 391 393 681 ICV_4 $T=853740 1092120 0 0 $X=853740 $Y=1091740
X499 1143 1 2 1146 404 405 681 ICV_4 $T=869860 1122360 0 0 $X=869860 $Y=1121980
X500 1169 1 2 1168 1166 1175 681 ICV_4 $T=891560 1102200 0 0 $X=891560 $Y=1101820
X501 413 1 2 415 416 418 681 ICV_4 $T=892800 1122360 0 0 $X=892800 $Y=1121980
X502 419 1 2 423 424 426 681 ICV_4 $T=902720 1122360 0 0 $X=902720 $Y=1121980
X503 1171 1 2 1179 1164 1174 681 ICV_4 $T=905820 1112280 1 0 $X=905820 $Y=1106860
X504 1188 1 2 1189 1190 1192 681 ICV_4 $T=924420 1122360 0 0 $X=924420 $Y=1121980
X505 1199 1 2 1201 451 454 681 ICV_4 $T=934340 1112280 1 0 $X=934340 $Y=1106860
X506 1205 1 2 1210 1187 1185 681 ICV_4 $T=941780 1122360 0 0 $X=941780 $Y=1121980
X507 455 1 2 458 459 465 681 ICV_4 $T=944260 1112280 1 0 $X=944260 $Y=1106860
X508 476 1 2 481 483 485 681 ICV_4 $T=964100 1122360 1 0 $X=964100 $Y=1116940
X509 488 1 2 491 473 494 681 ICV_4 $T=977120 1122360 0 0 $X=977120 $Y=1121980
X510 495 1 2 501 1240 1245 681 ICV_4 $T=987040 1112280 1 0 $X=987040 $Y=1106860
X511 1243 1 2 1244 498 1246 681 ICV_4 $T=992620 1092120 1 0 $X=992620 $Y=1086700
X512 1249 1 2 1248 510 515 681 ICV_4 $T=996960 1122360 1 0 $X=996960 $Y=1116940
X513 519 1 2 522 1265 1272 681 ICV_4 $T=1009360 1122360 0 0 $X=1009360 $Y=1121980
X514 1264 1 2 1261 523 1263 681 ICV_4 $T=1011220 1102200 0 0 $X=1011220 $Y=1101820
X515 1209 1 2 1226 529 532 681 ICV_4 $T=1020520 1122360 0 0 $X=1020520 $Y=1121980
X516 1283 1 2 1280 1285 1284 681 ICV_4 $T=1032920 1112280 1 0 $X=1032920 $Y=1106860
X517 1291 1 2 1294 1297 1298 681 ICV_4 $T=1048420 1112280 1 0 $X=1048420 $Y=1106860
X518 557 1 2 560 563 565 681 ICV_4 $T=1050280 1122360 0 0 $X=1050280 $Y=1121980
X519 1300 1 2 1301 571 577 681 ICV_4 $T=1058340 1112280 1 0 $X=1058340 $Y=1106860
X520 1307 1 2 1310 586 591 681 ICV_4 $T=1070740 1112280 1 0 $X=1070740 $Y=1106860
X521 601 1 2 1324 1326 1325 681 ICV_4 $T=1091200 1122360 1 0 $X=1091200 $Y=1116940
X522 608 1 2 610 611 615 681 ICV_4 $T=1091820 1122360 0 0 $X=1091820 $Y=1121980
X523 1330 1 2 1334 637 645 681 ICV_4 $T=1115380 1102200 1 0 $X=1115380 $Y=1096780
X524 755 1 2 757 58 62 681 ICV_5 $T=422220 1112280 0 0 $X=422220 $Y=1111900
X525 70 1 2 73 74 77 681 ICV_5 $T=436480 1122360 1 0 $X=436480 $Y=1116940
X526 105 1 2 108 110 117 681 ICV_5 $T=471200 1122360 0 0 $X=471200 $Y=1121980
X527 106 1 2 112 113 122 681 ICV_5 $T=474300 1122360 1 0 $X=474300 $Y=1116940
X528 120 1 2 125 128 134 681 ICV_5 $T=481740 1102200 1 0 $X=481740 $Y=1096780
X529 146 1 2 148 149 154 681 ICV_5 $T=505920 1122360 0 0 $X=505920 $Y=1121980
X530 173 1 2 176 178 183 681 ICV_5 $T=531960 1122360 0 0 $X=531960 $Y=1121980
X531 1091 1 2 1092 363 366 681 ICV_5 $T=809100 1112280 1 0 $X=809100 $Y=1106860
X532 1160 1 2 1162 410 412 681 ICV_5 $T=882880 1122360 0 0 $X=882880 $Y=1121980
X533 1296 1 2 1299 568 575 681 ICV_5 $T=1057100 1122360 1 0 $X=1057100 $Y=1116940
X534 574 1 2 579 580 584 681 ICV_5 $T=1065160 1122360 0 0 $X=1065160 $Y=1121980
X535 420 1 2 581 582 587 681 ICV_5 $T=1067020 1122360 1 0 $X=1067020 $Y=1116940
X536 585 1 2 589 592 597 681 ICV_5 $T=1075080 1122360 0 0 $X=1075080 $Y=1121980
X537 1230 1 2 1233 594 600 681 ICV_5 $T=1076940 1122360 1 0 $X=1076940 $Y=1116940
X538 1308 1 2 1322 629 633 681 ICV_5 $T=1106700 1122360 0 0 $X=1106700 $Y=1121980
X539 1329 1 2 1331 634 639 681 ICV_5 $T=1111660 1112280 1 0 $X=1111660 $Y=1106860
X540 724 39 2 1 720 36 MUX2 $T=389980 1092120 1 180 $X=385640 $Y=1091740
X541 728 39 2 1 719 37 MUX2 $T=389980 1102200 1 180 $X=385640 $Y=1101820
X542 730 41 2 1 721 37 MUX2 $T=390600 1102200 0 180 $X=386260 $Y=1096780
X543 733 41 2 1 723 40 MUX2 $T=394320 1102200 1 180 $X=389980 $Y=1101820
X544 738 39 2 1 736 40 MUX2 $T=399280 1102200 1 180 $X=394940 $Y=1101820
X545 51 49 2 1 734 36 MUX2 $T=406100 1092120 0 180 $X=401760 $Y=1086700
X546 742 49 2 1 740 37 MUX2 $T=406720 1102200 0 180 $X=402380 $Y=1096780
X547 748 49 2 1 741 747 MUX2 $T=416640 1102200 0 180 $X=412300 $Y=1096780
X548 751 49 2 1 743 53 MUX2 $T=418500 1092120 0 180 $X=414160 $Y=1086700
X549 758 41 2 1 750 57 MUX2 $T=427180 1102200 1 180 $X=422840 $Y=1101820
X550 757 39 2 1 761 66 MUX2 $T=432140 1102200 0 0 $X=432140 $Y=1101820
X551 764 41 2 1 762 66 MUX2 $T=439580 1092120 1 180 $X=435240 $Y=1091740
X552 763 39 2 1 766 765 MUX2 $T=437100 1102200 0 0 $X=437100 $Y=1101820
X553 770 81 2 1 768 765 MUX2 $T=450120 1102200 1 180 $X=445780 $Y=1101820
X554 773 81 2 1 769 747 MUX2 $T=455080 1102200 1 180 $X=450740 $Y=1101820
X555 783 81 2 1 772 36 MUX2 $T=463760 1092120 0 180 $X=459420 $Y=1086700
X556 786 101 2 1 780 765 MUX2 $T=467480 1102200 1 180 $X=463140 $Y=1101820
X557 793 101 2 1 782 747 MUX2 $T=474920 1112280 1 0 $X=474920 $Y=1106860
X558 799 127 2 1 795 747 MUX2 $T=486080 1112280 0 180 $X=481740 $Y=1106860
X559 121 101 2 1 800 129 MUX2 $T=483600 1092120 1 0 $X=483600 $Y=1086700
X560 803 127 2 1 797 130 MUX2 $T=492280 1092120 0 180 $X=487940 $Y=1086700
X561 808 127 2 1 802 765 MUX2 $T=496620 1112280 0 180 $X=492280 $Y=1106860
X562 810 127 2 1 805 129 MUX2 $T=498480 1092120 0 180 $X=494140 $Y=1086700
X563 818 147 2 1 812 144 MUX2 $T=507780 1102200 1 180 $X=503440 $Y=1101820
X564 817 147 2 1 806 765 MUX2 $T=507780 1112280 0 180 $X=503440 $Y=1106860
X565 819 151 2 1 814 765 MUX2 $T=512740 1112280 1 180 $X=508400 $Y=1111900
X566 164 147 2 1 815 150 MUX2 $T=522040 1092120 0 180 $X=517700 $Y=1086700
X567 828 151 2 1 826 144 MUX2 $T=525760 1112280 0 180 $X=521420 $Y=1106860
X568 827 151 2 1 824 150 MUX2 $T=527000 1092120 1 180 $X=522660 $Y=1091740
X569 834 151 2 1 829 171 MUX2 $T=533820 1092120 1 180 $X=529480 $Y=1091740
X570 832 151 2 1 833 836 MUX2 $T=532580 1112280 1 0 $X=532580 $Y=1106860
X571 181 147 2 1 838 171 MUX2 $T=538780 1092120 1 0 $X=538780 $Y=1086700
X572 837 147 2 1 839 836 MUX2 $T=541260 1112280 1 0 $X=541260 $Y=1106860
X573 843 193 2 1 840 171 MUX2 $T=551800 1092120 1 180 $X=547460 $Y=1091740
X574 845 193 2 1 842 836 MUX2 $T=553660 1112280 0 180 $X=549320 $Y=1106860
X575 852 193 2 1 846 169 MUX2 $T=561720 1112280 0 180 $X=557380 $Y=1106860
X576 857 206 2 1 850 171 MUX2 $T=566680 1102200 0 180 $X=562340 $Y=1096780
X577 860 193 2 1 865 219 MUX2 $T=572260 1102200 0 0 $X=572260 $Y=1101820
X578 862 206 2 1 863 169 MUX2 $T=572880 1112280 1 0 $X=572880 $Y=1106860
X579 864 206 2 1 868 219 MUX2 $T=575360 1092120 0 0 $X=575360 $Y=1091740
X580 871 206 2 1 872 867 MUX2 $T=582800 1112280 0 0 $X=582800 $Y=1111900
X581 880 881 2 1 875 169 MUX2 $T=597060 1112280 0 180 $X=592720 $Y=1106860
X582 873 228 2 1 232 189 MUX2 $T=593340 1092120 1 0 $X=593340 $Y=1086700
X583 884 237 2 1 877 169 MUX2 $T=603880 1112280 0 180 $X=599540 $Y=1106860
X584 890 240 2 1 882 885 MUX2 $T=610080 1092120 1 180 $X=605740 $Y=1091740
X585 891 881 2 1 878 885 MUX2 $T=610700 1102200 1 180 $X=606360 $Y=1101820
X586 894 237 2 1 887 885 MUX2 $T=611940 1112280 1 180 $X=607600 $Y=1111900
X587 907 237 2 1 900 867 MUX2 $T=619380 1112280 0 180 $X=615040 $Y=1106860
X588 912 881 2 1 910 867 MUX2 $T=628680 1102200 1 180 $X=624340 $Y=1101820
X589 911 228 2 1 914 867 MUX2 $T=624960 1092120 0 0 $X=624960 $Y=1091740
X590 870 240 2 1 908 867 MUX2 $T=633020 1102200 1 180 $X=628680 $Y=1101820
X591 918 240 2 1 916 219 MUX2 $T=637360 1102200 0 180 $X=633020 $Y=1096780
X592 259 228 2 1 256 257 MUX2 $T=637980 1092120 0 180 $X=633640 $Y=1086700
X593 921 240 2 1 917 257 MUX2 $T=642320 1102200 0 180 $X=637980 $Y=1096780
X594 923 237 2 1 913 929 MUX2 $T=642940 1112280 0 0 $X=642940 $Y=1111900
X595 934 881 2 1 922 929 MUX2 $T=651620 1112280 1 180 $X=647280 $Y=1111900
X596 933 881 2 1 927 267 MUX2 $T=652240 1102200 0 180 $X=647900 $Y=1096780
X597 936 881 2 1 939 257 MUX2 $T=652240 1112280 0 0 $X=652240 $Y=1111900
X598 273 228 2 1 275 267 MUX2 $T=652860 1092120 1 0 $X=652860 $Y=1086700
X599 946 237 2 1 948 944 MUX2 $T=660920 1112280 1 0 $X=660920 $Y=1106860
X600 947 237 2 1 949 267 MUX2 $T=666500 1102200 1 0 $X=666500 $Y=1096780
X601 954 283 2 1 956 929 MUX2 $T=672700 1112280 0 0 $X=672700 $Y=1111900
X602 957 289 2 1 951 929 MUX2 $T=681380 1112280 1 180 $X=677040 $Y=1111900
X603 966 296 2 1 963 929 MUX2 $T=688820 1102200 0 180 $X=684480 $Y=1096780
X604 969 298 2 1 967 929 MUX2 $T=692540 1112280 0 180 $X=688200 $Y=1106860
X605 970 298 2 1 973 971 MUX2 $T=693160 1112280 1 0 $X=693160 $Y=1106860
X606 975 289 2 1 964 971 MUX2 $T=699360 1112280 1 180 $X=695020 $Y=1111900
X607 981 298 2 1 984 982 MUX2 $T=703080 1112280 1 0 $X=703080 $Y=1106860
X608 986 289 2 1 978 982 MUX2 $T=708040 1122360 0 180 $X=703700 $Y=1116940
X609 990 296 2 1 979 267 MUX2 $T=711760 1092120 1 180 $X=707420 $Y=1091740
X610 997 289 2 1 1000 944 MUX2 $T=716100 1112280 0 0 $X=716100 $Y=1111900
X611 998 298 2 1 999 944 MUX2 $T=716720 1112280 1 0 $X=716720 $Y=1106860
X612 1006 283 2 1 1013 944 MUX2 $T=724780 1112280 0 0 $X=724780 $Y=1111900
X613 1017 283 2 1 1005 992 MUX2 $T=732840 1092120 1 180 $X=728500 $Y=1091740
X614 1010 296 2 1 1019 992 MUX2 $T=732220 1102200 1 0 $X=732220 $Y=1096780
X615 1018 296 2 1 1020 982 MUX2 $T=734080 1112280 1 0 $X=734080 $Y=1106860
X616 1021 283 2 1 1022 982 MUX2 $T=738420 1112280 1 0 $X=738420 $Y=1106860
X617 1015 316 2 1 1027 321 MUX2 $T=740900 1092120 1 0 $X=740900 $Y=1086700
X618 1023 296 2 1 1025 1028 MUX2 $T=742760 1112280 0 0 $X=742760 $Y=1111900
X619 1032 329 2 1 1024 1029 MUX2 $T=757640 1112280 1 180 $X=753300 $Y=1111900
X620 1036 329 2 1 1031 992 MUX2 $T=758880 1092120 1 180 $X=754540 $Y=1091740
X621 1041 329 2 1 1034 1028 MUX2 $T=763220 1112280 1 180 $X=758880 $Y=1111900
X622 1043 329 2 1 1033 294 MUX2 $T=766320 1092120 1 180 $X=761980 $Y=1091740
X623 1047 333 2 1 1038 1029 MUX2 $T=768800 1112280 1 180 $X=764460 $Y=1111900
X624 1048 333 2 1 1051 992 MUX2 $T=768800 1092120 0 0 $X=768800 $Y=1091740
X625 1055 333 2 1 1050 1028 MUX2 $T=773760 1112280 1 180 $X=769420 $Y=1111900
X626 1054 333 2 1 1049 1039 MUX2 $T=774380 1102200 1 180 $X=770040 $Y=1101820
X627 1065 343 2 1 1059 1039 MUX2 $T=786160 1092120 0 180 $X=781820 $Y=1086700
X628 1066 343 2 1 1062 992 MUX2 $T=786160 1102200 0 180 $X=781820 $Y=1096780
X629 1068 343 2 1 1064 1029 MUX2 $T=786780 1112280 1 180 $X=782440 $Y=1111900
X630 1079 343 2 1 1080 1028 MUX2 $T=794220 1112280 0 0 $X=794220 $Y=1111900
X631 1085 356 2 1 1082 352 MUX2 $T=804140 1092120 1 180 $X=799800 $Y=1091740
X632 1088 357 2 1 1083 1039 MUX2 $T=805380 1112280 1 180 $X=801040 $Y=1111900
X633 1092 356 2 1 1084 1029 MUX2 $T=809720 1112280 1 180 $X=805380 $Y=1111900
X634 362 356 2 1 1086 1039 MUX2 $T=813440 1092120 1 180 $X=809100 $Y=1091740
X635 1097 356 2 1 1100 369 MUX2 $T=817160 1092120 0 0 $X=817160 $Y=1091740
X636 1104 357 2 1 1095 1029 MUX2 $T=823360 1112280 1 180 $X=819020 $Y=1111900
X637 1102 357 2 1 1106 352 MUX2 $T=821500 1092120 0 0 $X=821500 $Y=1091740
X638 1105 357 2 1 1107 1028 MUX2 $T=823360 1112280 0 0 $X=823360 $Y=1111900
X639 1103 356 2 1 1113 1114 MUX2 $T=828320 1112280 1 0 $X=828320 $Y=1106860
X640 1110 374 2 1 1108 369 MUX2 $T=835760 1102200 0 180 $X=831420 $Y=1096780
X641 1116 374 2 1 1111 371 MUX2 $T=840100 1112280 0 180 $X=835760 $Y=1106860
X642 1115 374 2 1 1120 381 MUX2 $T=840100 1112280 1 0 $X=840100 $Y=1106860
X643 1124 383 2 1 1121 381 MUX2 $T=848780 1102200 1 180 $X=844440 $Y=1101820
X644 1125 383 2 1 1119 371 MUX2 $T=848780 1112280 1 180 $X=844440 $Y=1111900
X645 1131 374 2 1 1134 1114 MUX2 $T=853120 1112280 1 0 $X=853120 $Y=1106860
X646 1137 383 2 1 1139 1114 MUX2 $T=862420 1112280 0 180 $X=858080 $Y=1106860
X647 1146 399 2 1 1133 371 MUX2 $T=868000 1112280 0 180 $X=863660 $Y=1106860
X648 402 399 2 1 1155 369 MUX2 $T=872340 1092120 1 0 $X=872340 $Y=1086700
X649 1152 399 2 1 1149 1114 MUX2 $T=878540 1112280 1 180 $X=874200 $Y=1111900
X650 1154 399 2 1 1157 381 MUX2 $T=875440 1102200 0 0 $X=875440 $Y=1101820
X651 1128 406 2 1 1156 369 MUX2 $T=882260 1092120 0 180 $X=877920 $Y=1086700
X652 1162 406 2 1 1158 1114 MUX2 $T=883500 1112280 1 180 $X=879160 $Y=1111900
X653 1168 406 2 1 1163 381 MUX2 $T=888460 1112280 0 180 $X=884120 $Y=1106860
X654 1167 406 2 1 1170 371 MUX2 $T=887220 1102200 0 0 $X=887220 $Y=1101820
X655 1173 414 2 1 1172 1114 MUX2 $T=896520 1112280 0 180 $X=892180 $Y=1106860
X656 1174 414 2 1 1177 417 MUX2 $T=896520 1092120 0 0 $X=896520 $Y=1091740
X657 1175 414 2 1 1178 371 MUX2 $T=897140 1112280 1 0 $X=897140 $Y=1106860
X658 1179 414 2 1 1180 381 MUX2 $T=901480 1112280 1 0 $X=901480 $Y=1106860
X659 1185 433 2 1 1183 428 MUX2 $T=917600 1112280 1 180 $X=913260 $Y=1111900
X660 435 436 2 1 1184 428 MUX2 $T=920080 1092120 1 180 $X=915740 $Y=1091740
X661 1189 433 2 1 1181 442 MUX2 $T=924420 1102200 0 0 $X=924420 $Y=1101820
X662 443 436 2 1 1196 442 MUX2 $T=929380 1102200 1 0 $X=929380 $Y=1096780
X663 1192 436 2 1 1200 1197 MUX2 $T=929380 1112280 0 0 $X=929380 $Y=1111900
X664 1194 433 2 1 1191 1197 MUX2 $T=931240 1102200 0 0 $X=931240 $Y=1101820
X665 1201 433 2 1 1207 1204 MUX2 $T=934960 1102200 1 0 $X=934960 $Y=1096780
X666 1210 436 2 1 1202 1204 MUX2 $T=942400 1102200 1 180 $X=938060 $Y=1101820
X667 1216 436 2 1 1203 463 MUX2 $T=949220 1112280 0 0 $X=949220 $Y=1111900
X668 1223 469 2 1 1215 1204 MUX2 $T=959760 1102200 0 180 $X=955420 $Y=1096780
X669 1224 469 2 1 1217 428 MUX2 $T=959760 1112280 1 180 $X=955420 $Y=1111900
X670 1226 474 2 1 1220 1204 MUX2 $T=964100 1102200 0 180 $X=959760 $Y=1096780
X671 1231 469 2 1 1225 475 MUX2 $T=968440 1102200 0 180 $X=964100 $Y=1096780
X672 1227 474 2 1 1232 428 MUX2 $T=964720 1112280 0 0 $X=964720 $Y=1111900
X673 480 474 2 1 1234 475 MUX2 $T=968440 1102200 1 0 $X=968440 $Y=1096780
X674 484 474 2 1 1235 463 MUX2 $T=970300 1092120 0 0 $X=970300 $Y=1091740
X675 1233 469 2 1 1236 463 MUX2 $T=970300 1112280 0 0 $X=970300 $Y=1111900
X676 1245 503 2 1 1237 1197 MUX2 $T=992620 1112280 1 180 $X=988280 $Y=1111900
X677 1244 503 2 1 1241 1204 MUX2 $T=993240 1102200 0 180 $X=988900 $Y=1096780
X678 1246 504 2 1 1238 500 MUX2 $T=995720 1092120 1 180 $X=991380 $Y=1091740
X679 1248 506 2 1 1242 1197 MUX2 $T=997580 1112280 1 180 $X=993240 $Y=1111900
X680 1253 506 2 1 1247 1204 MUX2 $T=1000060 1102200 0 180 $X=995720 $Y=1096780
X681 1261 506 2 1 1250 428 MUX2 $T=1006880 1112280 0 180 $X=1002540 $Y=1106860
X682 1263 504 2 1 1268 520 MUX2 $T=1007500 1092120 1 0 $X=1007500 $Y=1086700
X683 1267 506 2 1 1271 475 MUX2 $T=1011220 1102200 1 0 $X=1011220 $Y=1096780
X684 1273 503 2 1 1266 521 MUX2 $T=1018040 1112280 1 180 $X=1013700 $Y=1111900
X685 1272 503 2 1 1270 475 MUX2 $T=1015560 1102200 1 0 $X=1015560 $Y=1096780
X686 1276 531 2 1 1274 521 MUX2 $T=1027960 1112280 1 180 $X=1023620 $Y=1111900
X687 1280 531 2 1 1275 500 MUX2 $T=1031680 1092120 1 180 $X=1027340 $Y=1091740
X688 1282 534 2 1 1278 521 MUX2 $T=1032920 1112280 0 180 $X=1028580 $Y=1106860
X689 1284 534 2 1 1281 535 MUX2 $T=1036640 1092120 1 180 $X=1032300 $Y=1091740
X690 540 541 2 1 536 535 MUX2 $T=1038500 1092120 0 180 $X=1034160 $Y=1086700
X691 1294 531 2 1 1288 553 MUX2 $T=1050900 1112280 1 180 $X=1046560 $Y=1111900
X692 554 541 2 1 1293 558 MUX2 $T=1047180 1092120 1 0 $X=1047180 $Y=1086700
X693 1298 531 2 1 1289 1292 MUX2 $T=1054620 1102200 0 180 $X=1050280 $Y=1096780
X694 1295 559 2 1 561 535 MUX2 $T=1051520 1092120 1 0 $X=1051520 $Y=1086700
X695 564 559 2 1 1302 558 MUX2 $T=1055860 1092120 1 0 $X=1055860 $Y=1086700
X696 1299 534 2 1 1303 553 MUX2 $T=1055860 1112280 0 0 $X=1055860 $Y=1111900
X697 1301 534 2 1 1304 1292 MUX2 $T=1058340 1102200 1 0 $X=1058340 $Y=1096780
X698 1310 593 2 1 1312 567 MUX2 $T=1083140 1092120 1 180 $X=1078800 $Y=1091740
X699 1317 599 2 1 1314 567 MUX2 $T=1087480 1092120 1 180 $X=1083140 $Y=1091740
X700 1319 605 2 1 1313 567 MUX2 $T=1090580 1112280 0 180 $X=1086240 $Y=1106860
X701 1322 609 2 1 1315 567 MUX2 $T=1094920 1112280 0 180 $X=1090580 $Y=1106860
X702 1324 609 2 1 1320 607 MUX2 $T=1096160 1092120 0 180 $X=1091820 $Y=1086700
X703 1325 599 2 1 1321 607 MUX2 $T=1096780 1092120 1 180 $X=1092440 $Y=1091740
X704 1327 605 2 1 1323 607 MUX2 $T=1099880 1112280 0 180 $X=1095540 $Y=1106860
X705 1331 605 2 1 1335 627 MUX2 $T=1107320 1112280 1 0 $X=1107320 $Y=1106860
X706 1333 599 2 1 1337 630 MUX2 $T=1110420 1092120 1 0 $X=1110420 $Y=1086700
X707 1334 599 2 1 1336 627 MUX2 $T=1111040 1102200 1 0 $X=1111040 $Y=1096780
X708 714 712 715 709 1 710 2 AOI22S $T=354640 1102200 1 180 $X=350920 $Y=1101820
X709 46 42 735 725 1 726 2 AOI22S $T=394940 1102200 0 180 $X=391220 $Y=1096780
X710 46 42 737 729 1 727 2 AOI22S $T=399280 1102200 0 180 $X=395560 $Y=1096780
X711 46 60 753 759 1 756 2 AOI22S $T=427800 1102200 0 0 $X=427800 $Y=1101820
X712 46 60 65 755 1 760 2 AOI22S $T=434620 1092120 0 180 $X=430900 $Y=1086700
X713 822 821 157 816 1 820 2 AOI22S $T=516460 1112280 0 180 $X=512740 $Y=1106860
X714 822 821 161 813 1 825 2 AOI22S $T=520800 1112280 0 180 $X=517080 $Y=1106860
X715 822 821 159 155 1 823 2 AOI22S $T=519560 1102200 1 0 $X=519560 $Y=1096780
X716 179 175 177 174 1 835 2 AOI22S $T=538160 1092120 1 180 $X=534440 $Y=1091740
X717 822 821 180 830 1 831 2 AOI22S $T=537540 1112280 1 0 $X=537540 $Y=1106860
X718 822 849 200 848 1 851 2 AOI22S $T=558620 1102200 1 0 $X=558620 $Y=1096780
X719 179 821 204 844 1 853 2 AOI22S $T=565440 1112280 0 180 $X=561720 $Y=1106860
X720 179 821 856 855 1 854 2 AOI22S $T=566680 1112280 1 0 $X=566680 $Y=1106860
X721 822 849 858 859 1 861 2 AOI22S $T=568540 1102200 1 0 $X=568540 $Y=1096780
X722 337 335 1056 1042 1 1026 2 AOI22S $T=777480 1092120 1 180 $X=773760 $Y=1091740
X723 337 335 1057 1053 1 1040 2 AOI22S $T=778100 1112280 1 180 $X=774380 $Y=1111900
X724 337 335 1058 1052 1 1044 2 AOI22S $T=778720 1102200 1 180 $X=775000 $Y=1101820
X725 337 335 1061 1046 1 1035 2 AOI22S $T=781820 1112280 1 180 $X=778100 $Y=1111900
X726 359 1090 1069 1089 1 1087 2 AOI22S $T=808480 1102200 0 180 $X=804760 $Y=1096780
X727 359 1090 1077 1093 1 360 2 AOI22S $T=808480 1102200 1 0 $X=808480 $Y=1096780
X728 359 1090 1072 1094 1 1091 2 AOI22S $T=810340 1112280 0 0 $X=810340 $Y=1111900
X729 359 1090 1081 1096 1 1098 2 AOI22S $T=814680 1112280 0 0 $X=814680 $Y=1111900
X730 1127 385 1130 1112 1 1118 2 AOI22S $T=852500 1102200 1 180 $X=848780 $Y=1101820
X731 1127 385 1126 1117 1 1122 2 AOI22S $T=853120 1112280 0 180 $X=849400 $Y=1106860
X732 386 385 1141 1132 1 1129 2 AOI22S $T=859940 1102200 0 0 $X=859940 $Y=1101820
X733 408 407 1153 1160 1 1159 2 AOI22S $T=883500 1102200 1 180 $X=879780 $Y=1101820
X734 408 407 1147 1123 1 1164 2 AOI22S $T=882260 1092120 1 0 $X=882260 $Y=1086700
X735 408 407 1140 1161 1 1166 2 AOI22S $T=883500 1102200 1 0 $X=883500 $Y=1096780
X736 408 407 1136 1169 1 1171 2 AOI22S $T=888460 1112280 1 0 $X=888460 $Y=1106860
X737 438 434 437 432 1 1187 2 AOI22S $T=922560 1092120 0 180 $X=918840 $Y=1086700
X738 438 434 441 439 1 1188 2 AOI22S $T=926280 1092120 0 180 $X=922560 $Y=1086700
X739 438 434 1195 1190 1 1186 2 AOI22S $T=930620 1092120 0 180 $X=926900 $Y=1086700
X740 438 434 448 1205 1 1199 2 AOI22S $T=936820 1092120 1 0 $X=936820 $Y=1086700
X741 1213 434 456 1212 1 453 2 AOI22S $T=946740 1092120 0 180 $X=943020 $Y=1086700
X742 1213 1218 461 1219 1 1221 2 AOI22S $T=952320 1092120 0 0 $X=952320 $Y=1091740
X743 1213 1218 468 1222 1 1209 2 AOI22S $T=957900 1092120 0 0 $X=957900 $Y=1091740
X744 1213 1218 471 1228 1 478 2 AOI22S $T=962240 1092120 0 0 $X=962240 $Y=1091740
X745 1213 1218 479 1230 1 482 2 AOI22S $T=965960 1092120 0 0 $X=965960 $Y=1091740
X746 1257 508 1256 1240 1 1249 2 AOI22S $T=1002540 1112280 0 180 $X=998820 $Y=1106860
X747 1257 508 1255 1243 1 1254 2 AOI22S $T=1004400 1102200 0 180 $X=1000680 $Y=1096780
X748 1257 508 516 1269 1 1264 2 AOI22S $T=1006880 1112280 1 0 $X=1006880 $Y=1106860
X749 1257 508 517 1265 1 1262 2 AOI22S $T=1007500 1102200 1 0 $X=1007500 $Y=1096780
X750 528 530 526 1279 1 1277 2 AOI22S $T=1025480 1102200 0 0 $X=1025480 $Y=1101820
X751 528 530 1252 1285 1 1283 2 AOI22S $T=1036640 1092120 0 0 $X=1036640 $Y=1091740
X752 542 543 1251 547 1 546 2 AOI22S $T=1039120 1092120 1 0 $X=1039120 $Y=1086700
X753 542 543 1259 549 1 552 2 AOI22S $T=1043460 1092120 1 0 $X=1043460 $Y=1086700
X754 528 1287 1258 1296 1 1291 2 AOI22S $T=1051520 1112280 0 0 $X=1051520 $Y=1111900
X755 528 1287 562 1300 1 1297 2 AOI22S $T=1054620 1102200 1 0 $X=1054620 $Y=1096780
X756 528 1287 1305 1307 1 1308 2 AOI22S $T=1065160 1102200 1 0 $X=1065160 $Y=1096780
X757 606 604 1306 1318 1 1316 2 AOI22S $T=1091820 1092120 1 180 $X=1088100 $Y=1091740
X758 606 604 612 1328 1 1326 2 AOI22S $T=1097400 1092120 0 0 $X=1097400 $Y=1091740
X759 606 604 617 1329 1 1330 2 AOI22S $T=1101740 1092120 0 0 $X=1101740 $Y=1091740
X760 606 604 623 624 1 1332 2 AOI22S $T=1106700 1092120 0 0 $X=1106700 $Y=1091740
X761 509 1255 1252 1251 2 1 505 AN4S $T=1001300 1092120 1 180 $X=996340 $Y=1091740
X762 511 1256 1258 1259 2 1 1198 AN4S $T=1002540 1092120 1 0 $X=1002540 $Y=1086700
X763 576 1306 1305 573 2 1 570 AN4S $T=1068260 1092120 0 180 $X=1063300 $Y=1086700
X764 5 2 1 6 BUF1 $T=282720 1092120 1 0 $X=282720 $Y=1086700
X765 55 2 1 29 BUF1 $T=363320 1122360 1 180 $X=360840 $Y=1121980
X766 30 2 1 694 BUF1 $T=367040 1112280 0 180 $X=364560 $Y=1106860
X767 53 2 1 57 BUF1 $T=440820 1092120 1 0 $X=440820 $Y=1086700
X768 111 2 1 788 BUF1 $T=475540 1092120 1 180 $X=473060 $Y=1091740
X769 114 2 1 790 BUF1 $T=479260 1092120 1 0 $X=479260 $Y=1086700
X770 747 2 1 135 BUF1 $T=488560 1112280 1 0 $X=488560 $Y=1106860
X771 150 2 1 130 BUF1 $T=512740 1092120 0 180 $X=510260 $Y=1086700
X772 30 2 1 170 BUF1 $T=527620 1102200 1 0 $X=527620 $Y=1096780
X773 150 2 1 189 BUF1 $T=543740 1092120 0 0 $X=543740 $Y=1091740
X774 30 2 1 841 BUF1 $T=545600 1112280 1 0 $X=545600 $Y=1106860
X775 175 2 1 849 BUF1 $T=556140 1092120 0 0 $X=556140 $Y=1091740
X776 849 2 1 821 BUF1 $T=570400 1112280 1 0 $X=570400 $Y=1106860
X777 257 2 1 944 BUF1 $T=657820 1112280 1 0 $X=657820 $Y=1106860
X778 317 2 1 982 BUF1 $T=736560 1092120 0 0 $X=736560 $Y=1091740
X779 944 2 1 1028 BUF1 $T=747720 1112280 0 0 $X=747720 $Y=1111900
X780 294 2 1 1039 BUF1 $T=758880 1092120 0 0 $X=758880 $Y=1091740
X781 992 2 1 352 BUF1 $T=792980 1092120 0 0 $X=792980 $Y=1091740
X782 365 2 1 1090 BUF1 $T=816540 1092120 1 180 $X=814060 $Y=1091740
X783 317 2 1 371 BUF1 $T=828320 1102200 1 0 $X=828320 $Y=1096780
X784 1028 2 1 1114 BUF1 $T=833280 1112280 1 0 $X=833280 $Y=1106860
X785 381 2 1 442 BUF1 $T=930000 1112280 1 0 $X=930000 $Y=1106860
X786 447 2 1 1213 BUF1 $T=949840 1092120 0 0 $X=949840 $Y=1091740
X787 514 2 1 1257 BUF1 $T=1006880 1102200 0 180 $X=1004400 $Y=1096780
X788 500 2 1 535 BUF1 $T=1030440 1092120 1 0 $X=1030440 $Y=1086700
X789 475 2 1 551 BUF1 $T=1046560 1102200 1 0 $X=1046560 $Y=1096780
X790 567 2 1 558 BUF1 $T=1060200 1092120 1 0 $X=1060200 $Y=1086700
X791 553 2 1 567 BUF1 $T=1062680 1102200 1 0 $X=1062680 $Y=1096780
X792 1030 1 2 1032 BUF1CK $T=752680 1112280 1 0 $X=752680 $Y=1106860
X793 1037 1 2 1036 BUF1CK $T=761360 1092120 1 0 $X=761360 $Y=1086700
X794 1101 1 2 1103 BUF1CK $T=820260 1112280 1 0 $X=820260 $Y=1106860
X795 1176 1 2 1173 BUF1CK $T=901480 1102200 0 0 $X=901480 $Y=1101820
X796 1193 1 2 1194 BUF1CK $T=935580 1102200 0 0 $X=935580 $Y=1101820
X797 1206 1 2 1208 BUF1CK $T=939300 1122360 0 0 $X=939300 $Y=1121980
X798 1229 1 2 1227 BUF1CK $T=972160 1112280 1 0 $X=972160 $Y=1106860
X799 530 1 2 1287 BUF1CK $T=1042840 1102200 1 0 $X=1042840 $Y=1096780
X800 1214 434 1 2 INV2 $T=946740 1092120 1 0 $X=946740 $Y=1086700
X801 518 513 1 2 INV2 $T=1008120 1122360 1 180 $X=1006260 $Y=1121980
X802 1109 1110 1 2 BUF2 $T=827700 1122360 1 0 $X=827700 $Y=1116940
X803 375 1109 1 2 BUF2 $T=838860 1092120 1 0 $X=838860 $Y=1086700
X804 1212 1206 1 2 BUF2 $T=949220 1122360 1 0 $X=949220 $Y=1116940
X805 15 1 689 693 2 17 ND3 $T=325500 1102200 1 0 $X=325500 $Y=1096780
X806 24 1 709 708 2 22 ND3 $T=347200 1092120 0 180 $X=344720 $Y=1086700
X807 731 1 43 732 2 735 ND3 $T=393080 1092120 1 0 $X=393080 $Y=1086700
X808 745 1 50 744 2 737 ND3 $T=409820 1102200 0 180 $X=407340 $Y=1096780
X809 749 1 54 754 2 753 ND3 $T=417880 1102200 0 0 $X=417880 $Y=1101820
X810 856 1 213 217 2 798 ND3 $T=572260 1092120 1 0 $X=572260 $Y=1086700
X811 858 1 214 210 2 779 ND3 $T=572260 1092120 0 0 $X=572260 $Y=1091740
X812 1070 1 1069 345 2 1056 ND3 $T=789880 1102200 0 180 $X=787400 $Y=1096780
X813 1071 1 1072 348 2 1061 ND3 $T=789260 1112280 0 0 $X=789260 $Y=1111900
X814 1076 1 1077 350 2 1058 ND3 $T=792980 1102200 1 0 $X=792980 $Y=1096780
X815 1078 1 1081 354 2 1057 ND3 $T=797940 1112280 1 0 $X=797940 $Y=1106860
X816 1135 1 1130 389 2 1136 ND3 $T=854980 1102200 0 0 $X=854980 $Y=1101820
X817 1138 1 1126 392 2 1140 ND3 $T=857460 1102200 0 0 $X=857460 $Y=1101820
X818 1150 1 398 397 2 1147 ND3 $T=867380 1092120 1 0 $X=867380 $Y=1086700
X819 1151 1 1141 403 2 1153 ND3 $T=872340 1112280 1 0 $X=872340 $Y=1106860
X820 444 1 1195 445 2 1198 ND3 $T=931240 1092120 1 0 $X=931240 $Y=1086700
X821 13 691 695 2 1 ND2S $T=318680 1092120 0 0 $X=318680 $Y=1091740
X822 689 692 15 2 1 ND2S $T=322400 1102200 1 0 $X=322400 $Y=1096780
X823 17 698 15 2 1 ND2S $T=329840 1102200 0 180 $X=327980 $Y=1096780
X824 705 704 697 2 1 ND2S $T=340380 1092120 1 180 $X=338520 $Y=1091740
X825 27 26 25 2 1 ND2S $T=350920 1092120 0 180 $X=349060 $Y=1086700
X826 44 45 47 2 1 ND2S $T=395560 1092120 1 0 $X=395560 $Y=1086700
X827 44 731 739 2 1 ND2S $T=400520 1102200 1 0 $X=400520 $Y=1096780
X828 44 745 746 2 1 ND2S $T=409820 1102200 1 0 $X=409820 $Y=1096780
X829 44 749 752 2 1 ND2S $T=416640 1102200 1 0 $X=416640 $Y=1096780
X830 346 1070 1063 2 1 ND2S $T=789260 1102200 1 180 $X=787400 $Y=1101820
X831 346 1071 1067 2 1 ND2S $T=789260 1112280 1 180 $X=787400 $Y=1111900
X832 346 1076 1074 2 1 ND2S $T=792360 1102200 0 180 $X=790500 $Y=1096780
X833 346 1078 1075 2 1 ND2S $T=793600 1112280 1 180 $X=791740 $Y=1111900
X834 401 1138 1143 2 1 ND2S $T=864280 1102200 0 0 $X=864280 $Y=1101820
X835 401 1135 1145 2 1 ND2S $T=869240 1102200 0 0 $X=869240 $Y=1101820
X836 401 1151 1148 2 1 ND2S $T=869240 1112280 1 0 $X=869240 $Y=1106860
X837 401 1150 400 2 1 ND2S $T=869860 1092120 1 0 $X=869860 $Y=1086700
X838 686 8 1 685 684 682 2 MOAI1S $T=300080 1092120 0 180 $X=296360 $Y=1086700
X839 690 693 1 692 691 687 2 MOAI1S $T=316200 1102200 0 180 $X=312480 $Y=1096780
X840 689 698 1 689 698 699 2 MOAI1S $T=329840 1102200 1 0 $X=329840 $Y=1096780
X841 713 711 1 713 711 716 2 MOAI1S $T=352160 1092120 0 0 $X=352160 $Y=1091740
X842 790 102 1 788 784 787 2 MOAI1S $T=471820 1092120 0 180 $X=468100 $Y=1086700
X843 790 785 1 788 775 778 2 MOAI1S $T=471820 1102200 1 180 $X=468100 $Y=1101820
X844 790 791 1 788 777 794 2 MOAI1S $T=471820 1102200 0 0 $X=471820 $Y=1101820
X845 790 109 1 111 792 796 2 MOAI1S $T=475540 1092120 1 0 $X=475540 $Y=1086700
X846 893 889 1 896 897 899 2 MOAI1S $T=610700 1102200 1 0 $X=610700 $Y=1096780
X847 893 879 1 896 888 245 2 MOAI1S $T=610700 1102200 0 0 $X=610700 $Y=1101820
X848 243 222 1 244 892 898 2 MOAI1S $T=611940 1092120 0 0 $X=611940 $Y=1091740
X849 243 901 1 244 905 904 2 MOAI1S $T=618140 1102200 1 0 $X=618140 $Y=1096780
X850 893 902 1 896 906 909 2 MOAI1S $T=618140 1102200 0 0 $X=618140 $Y=1101820
X851 243 264 1 250 925 926 2 MOAI1S $T=641080 1092120 1 0 $X=641080 $Y=1086700
X852 243 271 1 250 928 931 2 MOAI1S $T=652860 1092120 0 180 $X=649140 $Y=1086700
X853 893 937 1 272 932 269 2 MOAI1S $T=654720 1112280 0 180 $X=651000 $Y=1106860
X854 893 935 1 272 938 930 2 MOAI1S $T=652860 1102200 1 0 $X=652860 $Y=1096780
X855 893 941 1 272 945 943 2 MOAI1S $T=657820 1102200 1 0 $X=657820 $Y=1096780
X856 276 955 1 272 952 953 2 MOAI1S $T=675180 1092120 1 180 $X=671460 $Y=1091740
X857 295 959 1 293 962 961 2 MOAI1S $T=688200 1112280 0 180 $X=684480 $Y=1106860
X858 295 965 1 293 977 974 2 MOAI1S $T=698120 1112280 1 0 $X=698120 $Y=1106860
X859 295 980 1 293 987 988 2 MOAI1S $T=708040 1112280 1 0 $X=708040 $Y=1106860
X860 295 991 1 293 994 995 2 MOAI1S $T=712380 1112280 1 0 $X=712380 $Y=1106860
X861 312 1007 1 311 1004 1002 2 MOAI1S $T=727260 1112280 0 180 $X=723540 $Y=1106860
X862 312 1001 1 311 1008 976 2 MOAI1S $T=731600 1102200 0 180 $X=727880 $Y=1096780
X863 312 1011 1 311 1016 1012 2 MOAI1S $T=729740 1112280 1 0 $X=729740 $Y=1106860
X864 695 2 697 692 1 NR2 $T=322400 1092120 0 0 $X=322400 $Y=1091740
X865 706 2 20 708 1 NR2 $T=341620 1092120 1 0 $X=341620 $Y=1086700
X866 709 2 25 704 1 NR2 $T=347200 1092120 0 0 $X=347200 $Y=1091740
X867 707 2 710 704 1 NR2 $T=347200 1102200 0 0 $X=347200 $Y=1101820
X868 707 2 711 26 1 NR2 $T=349060 1092120 0 0 $X=349060 $Y=1091740
X869 778 2 779 754 1 NR2 $T=458800 1102200 0 0 $X=458800 $Y=1101820
X870 787 2 97 98 1 NR2 $T=468100 1092120 0 180 $X=466240 $Y=1086700
X871 794 2 115 744 1 NR2 $T=476780 1102200 0 0 $X=476780 $Y=1101820
X872 796 2 798 732 1 NR2 $T=481740 1092120 1 0 $X=481740 $Y=1086700
X873 898 2 249 899 1 NR2 $T=615040 1102200 1 0 $X=615040 $Y=1096780
X874 904 2 251 909 1 NR2 $T=620620 1092120 0 0 $X=620620 $Y=1091740
X875 926 2 268 930 1 NR2 $T=646660 1092120 1 0 $X=646660 $Y=1086700
X876 931 2 277 943 1 NR2 $T=657820 1092120 1 0 $X=657820 $Y=1086700
X877 961 2 291 953 1 NR2 $T=684480 1102200 0 180 $X=682620 $Y=1096780
X878 974 2 303 976 1 NR2 $T=698740 1102200 1 0 $X=698740 $Y=1096780
X879 995 2 309 1002 1 NR2 $T=721680 1112280 1 0 $X=721680 $Y=1106860
X880 988 2 313 1012 1 NR2 $T=727260 1112280 1 0 $X=727260 $Y=1106860
X881 3 4 1 2 INV12CK $T=220100 1122360 0 0 $X=220100 $Y=1121980
X882 4 38 1 2 INV12CK $T=393080 1092120 0 180 $X=383160 $Y=1086700
X883 705 21 2 1 706 OR2 $T=344100 1092120 1 180 $X=341620 $Y=1091740
X884 705 701 19 704 2 1 703 OA22 $T=341000 1102200 0 180 $X=336660 $Y=1096780
X885 13 697 1 2 701 AN2 $T=334180 1102200 1 0 $X=334180 $Y=1096780
X886 686 2 689 690 12 1 NR3 $T=308760 1102200 1 0 $X=308760 $Y=1096780
X887 686 9 1 684 2 OR2B1S $T=304420 1092120 0 180 $X=301320 $Y=1086700
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=15 FDC=0
X0 1 2 3 4 5 6 MUX2 $T=4340 0 0 0 $X=4340 $Y=-380
X1 7 8 9 10 4 11 3 AOI22S $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 DELB $T=0 0 0 0 $X=0 $Y=-380
X1 5 6 7 3 2 8 QDFFRBN $T=16740 0 1 180 $X=4960 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=15 FDC=0
X0 1 2 3 4 5 6 MUX2 $T=3720 0 0 0 $X=3720 $Y=-380
X1 7 8 9 10 4 11 3 AOI22S $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 DELB $T=0 0 1 180 $X=-4960 $Y=-380
X1 5 6 7 3 2 8 QDFFRBN $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 DELB $T=0 0 0 0 $X=0 $Y=-380
X1 5 6 7 3 2 8 QDFFRBN $T=4960 0 0 0 $X=4960 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 INV1S $T=0 0 0 0 $X=0 $Y=-380
X1 5 6 7 2 4 8 QDFFRBN $T=1240 0 0 0 $X=1240 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=15 FDC=0
X0 1 2 3 4 5 6 MUX2 $T=0 0 0 0 $X=0 $Y=-380
X1 7 8 9 10 4 11 3 AOI22S $T=-3720 0 0 0 $X=-3720 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=0
X0 1 2 3 4 BUF1S $T=4960 0 0 0 $X=4960 $Y=-380
X1 5 2 3 6 DELB $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 DELB $T=11780 0 0 0 $X=11780 $Y=-380
X1 5 6 7 3 2 8 QDFFRBN $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=0
X0 1 2 3 4 INV1S $T=0 0 0 0 $X=0 $Y=-380
X1 5 2 6 4 INV1S $T=1240 0 0 0 $X=1240 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=0
X0 1 2 3 4 INV1S $T=4960 0 0 0 $X=4960 $Y=-380
X1 5 4 2 6 DELB $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT INV6CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN4 I1 I2 I4 I3 O GND VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR3H O I3 I2 I1 VCC GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND2 I1 O I2 GND VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA112 A1 B1 C1 C2 VCC GND O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV8CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI112HS C2 C1 GND B1 O A1 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22HP A2 A1 VCC B1 O B2 GND
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22H A2 A1 VCC B1 O B2 GND
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND3P I1 O I2 I3 GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR2P I1 VCC I2 GND O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN4B1S I3 I2 I1 VCC B1 GND O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF3CK I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FA1S CO VCC A B CI GND S
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNR2HS I1 I2 O VCC GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA12 B2 B1 A1 GND VCC O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI22S B2 GND B1 A2 O A1 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO22 O A2 A1 VCC B1 B2 GND
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MUX3 B S0 A S1 VCC C GND O
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO12 B2 B1 A1 GND VCC O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI12HS B2 B1 VCC A1 GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN2B1S I1 VCC B1 O GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI12HS B2 B1 GND A1 VCC O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MAOI1 B1 B2 A1 A2 VCC GND O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR3B2S I1 B1 VCC O B2 GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MOAI1 B1 B2 GND A1 O A2 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540
+ 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560
+ 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580
+ 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640
+ 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660
+ 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680
+ 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700
+ 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720
+ 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740
+ 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760
+ 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780
+ 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800
+ 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820
+ 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840
+ 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860
+ 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880
+ 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900
+ 901 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920
+ 921 922 923 924 925 926 927 928 929 930 931 932 933 934 935 936 937 938 939 940
+ 941 942 943 944 945 946 947 948 949 950 951 952 953 954 955 956 957 958 959 960
+ 961 962 963 964 965 966 967 968 969 970 971 972 973 974 975 976 977 978 979 980
+ 981 982 983 984 985 986 987 988 989 990 991 992 993 994 995 996 997 998 999 1000
+ 1001 1002 1003 1004 1005 1006 1007 1008 1009 1010 1011 1012 1013 1014 1015 1016 1017 1018 1019 1020
+ 1021 1022 1023 1024 1025 1026 1027 1028 1029 1030 1031 1032 1033 1034 1035 1036 1037 1038 1039 1040
+ 1041 1042 1043 1044 1045 1046 1047 1048 1049 1050 1051 1052 1053 1054 1055 1056 1057 1058 1059 1060
+ 1061 1062 1063 1064 1065 1066 1067 1068 1069 1070 1071 1072 1073 1074 1075 1076 1077 1078 1079 1080
+ 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 1093 1094 1095 1096 1097 1098 1099 1100
+ 1101 1102 1103 1104 1105 1106 1107 1108 1109 1110 1111 1112 1113 1114 1115 1116 1117 1118 1119 1120
+ 1121 1122 1123 1124 1125 1126 1127 1128 1129 1130 1131 1132 1133 1134 1135 1136 1137 1138 1139 1140
+ 1141 1142 1143 1144 1145 1146 1147 1148 1149 1150 1151 1152 1153 1154 1155 1156 1157 1158 1159 1160
+ 1161 1162 1163 1164 1165 1166 1167 1168 1169 1170 1171 1172 1173 1174 1175 1176 1177 1178 1179 1180
+ 1181 1182 1183 1184 1185 1186 1187 1188 1189 1190 1191 1192 1193 1194 1195 1196 1197 1198 1199 1200
+ 1201 1202 1203 1204 1205 1206 1207 1208 1209 1210 1211 1212 1213 1214 1215 1216 1217 1218 1219 1220
+ 1221 1222 1223 1224 1225 1226 1227 1228 1229 1230 1231 1232 1233 1234 1235 1236 1237 1238 1239 1240
+ 1241 1242 1243 1244 1245 1246 1247 1248 1249 1250 1251 1252 1253 1254 1255 1256 1257 1258 1259 1260
+ 1261 1262 1263 1264 1265 1266 1267 1268 1269 1270 1271 1272 1273 1274 1275 1276 1277 1278 1279 1280
+ 1281 1282 1283 1284 1285 1286 1287 1288 1289 1291 1299
** N=6533 EP=1291 IP=34617 FDC=0
X0 1288 6532 6532 6532 1291 6532 1289 YA2GSD $T=1349740 983520 0 90 $X=1210240 $Y=986370
X1 1302 2 1327 1 INV1S $T=224440 1061880 1 0 $X=224440 $Y=1056460
X2 1301 2 1328 1 INV1S $T=225680 920760 1 0 $X=225680 $Y=915340
X3 1312 2 1343 1 INV1S $T=226300 930840 0 0 $X=226300 $Y=930460
X4 1351 2 1329 1 INV1S $T=227540 940920 1 180 $X=226300 $Y=940540
X5 1313 2 1344 1 INV1S $T=226300 951000 0 0 $X=226300 $Y=950620
X6 1303 2 1356 1 INV1S $T=228160 920760 0 0 $X=228160 $Y=920380
X7 1353 2 1352 1 INV1S $T=228160 971160 1 0 $X=228160 $Y=965740
X8 1347 2 1359 1 INV1S $T=228160 1051800 0 0 $X=228160 $Y=1051420
X9 1363 2 1379 1 INV1S $T=230020 920760 0 0 $X=230020 $Y=920380
X10 1385 2 1318 1 INV1S $T=233120 910680 0 180 $X=231880 $Y=905260
X11 1366 2 1426 1 INV1S $T=233740 951000 1 0 $X=233740 $Y=945580
X12 1348 2 1398 1 INV1S $T=233740 971160 0 0 $X=233740 $Y=970780
X13 1394 2 1406 1 INV1S $T=233740 1071960 1 0 $X=233740 $Y=1066540
X14 1409 2 1376 1 INV1S $T=236220 910680 0 180 $X=234980 $Y=905260
X15 1444 2 1404 1 INV1S $T=236840 920760 1 180 $X=235600 $Y=920380
X16 1357 2 1425 1 INV1S $T=235600 940920 1 0 $X=235600 $Y=935500
X17 1368 2 1412 1 INV1S $T=235600 1061880 0 0 $X=235600 $Y=1061500
X18 1440 2 1396 1 INV1S $T=239940 961080 0 180 $X=238700 $Y=955660
X19 1443 2 1449 1 INV1S $T=241180 1082040 1 0 $X=241180 $Y=1076620
X20 1471 2 1445 1 INV1S $T=245520 930840 1 180 $X=244280 $Y=930460
X21 1450 2 1455 1 INV1S $T=245520 940920 0 0 $X=245520 $Y=940540
X22 1486 2 1465 1 INV1S $T=247380 910680 1 180 $X=246140 $Y=910300
X23 1531 2 1480 1 INV1S $T=249240 961080 1 180 $X=248000 $Y=960700
X24 1485 2 1502 1 INV1S $T=248620 1082040 1 0 $X=248620 $Y=1076620
X25 1517 2 1476 1 INV1S $T=252340 971160 1 180 $X=251100 $Y=970780
X26 1529 2 1456 1 INV1S $T=254200 910680 1 180 $X=252960 $Y=910300
X27 1534 2 1501 1 INV1S $T=254200 1041720 1 180 $X=252960 $Y=1041340
X28 1555 2 1568 1 INV1S $T=257920 1051800 1 0 $X=257920 $Y=1046380
X29 1561 2 1569 1 INV1S $T=258540 1082040 1 0 $X=258540 $Y=1076620
X30 32 2 38 1 INV1S $T=259780 930840 0 0 $X=259780 $Y=930460
X31 1542 2 1574 1 INV1S $T=260400 920760 1 0 $X=260400 $Y=915340
X32 1581 2 1571 1 INV1S $T=261640 971160 0 180 $X=260400 $Y=965740
X33 1544 2 1591 1 INV1S $T=261020 1031640 1 0 $X=261020 $Y=1026220
X34 1586 2 1560 1 INV1S $T=262880 1021560 0 180 $X=261640 $Y=1016140
X35 1613 2 1578 1 INV1S $T=265360 1041720 0 180 $X=264120 $Y=1036300
X36 1612 2 29 1 INV1S $T=269080 1031640 0 180 $X=267840 $Y=1026220
X37 1620 2 1648 1 INV1S $T=267840 1061880 1 0 $X=267840 $Y=1056460
X38 1589 2 1636 1 INV1S $T=268460 930840 1 0 $X=268460 $Y=925420
X39 1550 2 50 1 INV1S $T=272180 910680 0 180 $X=270940 $Y=905260
X40 54 2 48 1 INV1S $T=272800 900600 1 180 $X=271560 $Y=900220
X41 1644 2 1643 1 INV1S $T=272800 1021560 0 180 $X=271560 $Y=1016140
X42 1549 2 1667 1 INV1S $T=272800 1071960 0 0 $X=272800 $Y=1071580
X43 1612 2 1677 1 INV1S $T=274040 1041720 1 0 $X=274040 $Y=1036300
X44 53 2 55 1 INV1S $T=274660 910680 1 0 $X=274660 $Y=905260
X45 1730 2 1685 1 INV1S $T=283340 961080 0 180 $X=282100 $Y=955660
X46 1731 2 1622 1 INV1S $T=283960 940920 1 180 $X=282720 $Y=940540
X47 62 2 1737 1 INV1S $T=286440 910680 1 180 $X=285200 $Y=910300
X48 1752 2 1817 1 INV1S $T=287060 1082040 1 0 $X=287060 $Y=1076620
X49 1509 2 1618 1 INV1S $T=288920 1001400 0 180 $X=287680 $Y=995980
X50 1744 2 1763 1 INV1S $T=288300 940920 1 0 $X=288300 $Y=935500
X51 1758 2 1774 1 INV1S $T=289540 1051800 0 0 $X=289540 $Y=1051420
X52 1784 2 1765 1 INV1S $T=292020 951000 1 180 $X=290780 $Y=950620
X53 1541 2 1657 1 INV1S $T=292640 1021560 1 0 $X=292640 $Y=1016140
X54 1785 2 1816 1 INV1S $T=295120 1031640 0 0 $X=295120 $Y=1031260
X55 59 2 1822 1 INV1S $T=295740 910680 1 0 $X=295740 $Y=905260
X56 68 2 1820 1 INV1S $T=295740 1021560 1 0 $X=295740 $Y=1016140
X57 1815 2 1809 1 INV1S $T=295740 1061880 0 0 $X=295740 $Y=1061500
X58 1762 2 65 1 INV1S $T=297600 930840 0 180 $X=296360 $Y=925420
X59 1812 2 1845 1 INV1S $T=298220 971160 1 0 $X=298220 $Y=965740
X60 1837 2 1846 1 INV1S $T=298220 1061880 0 0 $X=298220 $Y=1061500
X61 1853 2 1832 1 INV1S $T=300080 930840 1 180 $X=298840 $Y=930460
X62 1618 2 1854 1 INV1S $T=299460 1001400 1 0 $X=299460 $Y=995980
X63 1825 2 1857 1 INV1S $T=299460 1071960 1 0 $X=299460 $Y=1066540
X64 1854 2 1639 1 INV1S $T=300080 1011480 1 0 $X=300080 $Y=1006060
X65 1822 2 1813 1 INV1S $T=302560 920760 0 180 $X=301320 $Y=915340
X66 1674 2 1863 1 INV1S $T=301940 1031640 1 0 $X=301940 $Y=1026220
X67 79 2 1612 1 INV1S $T=304420 1031640 0 180 $X=303180 $Y=1026220
X68 1896 2 1716 1 INV1S $T=306900 1011480 0 180 $X=305660 $Y=1006060
X69 1894 2 1883 1 INV1S $T=306900 961080 1 0 $X=306900 $Y=955660
X70 1854 2 1903 1 INV1S $T=306900 1001400 1 0 $X=306900 $Y=995980
X71 1896 2 1910 1 INV1S $T=308140 1001400 0 0 $X=308140 $Y=1001020
X72 75 2 1896 1 INV1S $T=309380 1011480 0 180 $X=308140 $Y=1006060
X73 1944 2 83 1 INV1S $T=311240 981240 1 180 $X=310000 $Y=980860
X74 1930 2 1893 1 INV1S $T=311860 1051800 0 180 $X=310620 $Y=1046380
X75 1931 2 1918 1 INV1S $T=313720 961080 1 180 $X=312480 $Y=960700
X76 1940 2 1946 1 INV1S $T=313720 1071960 1 0 $X=313720 $Y=1066540
X77 111 2 1928 1 INV1S $T=319300 920760 1 180 $X=318060 $Y=920380
X78 1926 2 1965 1 INV1S $T=319300 1031640 1 180 $X=318060 $Y=1031260
X79 115 2 1953 1 INV1S $T=319920 1082040 1 180 $X=318680 $Y=1081660
X80 106 2 1911 1 INV1S $T=319300 910680 0 0 $X=319300 $Y=910300
X81 112 2 99 1 INV1S $T=321780 930840 0 180 $X=320540 $Y=925420
X82 1988 2 108 1 INV1S $T=323640 1021560 0 180 $X=322400 $Y=1016140
X83 1550 2 1974 1 INV1S $T=323020 920760 1 0 $X=323020 $Y=915340
X84 1989 2 74 1 INV1S $T=324260 991320 1 0 $X=324260 $Y=985900
X85 1906 2 1968 1 INV1S $T=326120 930840 0 0 $X=326120 $Y=930460
X86 2003 2 2014 1 INV1S $T=326740 940920 1 0 $X=326740 $Y=935500
X87 1997 2 92 1 INV1S $T=327360 991320 1 0 $X=327360 $Y=985900
X88 2026 2 2008 1 INV1S $T=329220 1061880 1 180 $X=327980 $Y=1061500
X89 2024 2 123 1 INV1S $T=329840 1021560 0 180 $X=328600 $Y=1016140
X90 2019 2 117 1 INV1S $T=331080 1082040 1 0 $X=331080 $Y=1076620
X91 2054 2 2030 1 INV1S $T=332940 1071960 1 180 $X=331700 $Y=1071580
X92 2038 2 2042 1 INV1S $T=333560 930840 1 180 $X=332320 $Y=930460
X93 2071 2 128 1 INV1S $T=337280 940920 0 180 $X=336040 $Y=935500
X94 2098 2 2081 1 INV1S $T=339140 1071960 0 180 $X=337900 $Y=1066540
X95 1822 2 146 1 INV1S $T=340380 900600 0 0 $X=340380 $Y=900220
X96 140 2 2115 1 INV1S $T=340380 1061880 1 0 $X=340380 $Y=1056460
X97 2111 2 2134 1 INV1S $T=340380 1071960 0 0 $X=340380 $Y=1071580
X98 2146 2 1849 1 INV1S $T=344720 1061880 0 180 $X=343480 $Y=1056460
X99 2153 2 2176 1 INV1S $T=347200 940920 0 0 $X=347200 $Y=940540
X100 159 2 2137 1 INV1S $T=348440 1082040 1 180 $X=347200 $Y=1081660
X101 161 2 155 1 INV1S $T=350300 1082040 0 180 $X=349060 $Y=1076620
X102 2157 2 2185 1 INV1S $T=350920 951000 0 0 $X=350920 $Y=950620
X103 2187 2 2196 1 INV1S $T=352160 940920 1 0 $X=352160 $Y=935500
X104 2159 2 2202 1 INV1S $T=353400 1021560 1 0 $X=353400 $Y=1016140
X105 2163 2 2129 1 INV1S $T=354640 1051800 0 180 $X=353400 $Y=1046380
X106 2210 2 2182 1 INV1S $T=355880 1021560 0 180 $X=354640 $Y=1016140
X107 2228 2 2212 1 INV1S $T=358980 951000 0 180 $X=357740 $Y=945580
X108 2225 2 2237 1 INV1S $T=358980 910680 0 0 $X=358980 $Y=910300
X109 2260 2 1669 1 INV1S $T=362700 1061880 0 180 $X=361460 $Y=1056460
X110 2240 2 2263 1 INV1S $T=364560 961080 1 0 $X=364560 $Y=955660
X111 2308 2 2245 1 INV1S $T=366420 910680 0 180 $X=365180 $Y=905260
X112 2266 2 2255 1 INV1S $T=366420 971160 1 180 $X=365180 $Y=970780
X113 2128 2 2204 1 INV1S $T=365180 1001400 1 0 $X=365180 $Y=995980
X114 162 2 2284 1 INV1S $T=368280 1001400 0 0 $X=368280 $Y=1001020
X115 2220 2 2194 1 INV1S $T=370140 1041720 1 180 $X=368900 $Y=1041340
X116 184 2 2275 1 INV1S $T=370760 1061880 0 0 $X=370760 $Y=1061500
X117 2279 2 2338 1 INV1S $T=374480 971160 1 0 $X=374480 $Y=965740
X118 2327 2 2358 1 INV1S $T=377580 951000 1 0 $X=377580 $Y=945580
X119 2331 2 2364 1 INV1S $T=377580 971160 1 0 $X=377580 $Y=965740
X120 2376 2 2345 1 INV1S $T=378820 981240 0 180 $X=377580 $Y=975820
X121 2377 2 2233 1 INV1S $T=380680 1001400 1 180 $X=379440 $Y=1001020
X122 2275 2 2373 1 INV1S $T=383160 1041720 1 180 $X=381920 $Y=1041340
X123 2246 2 2403 1 INV1S $T=385020 940920 1 0 $X=385020 $Y=935500
X124 2401 2 2407 1 INV1S $T=385640 971160 0 0 $X=385640 $Y=970780
X125 2377 2 2394 1 INV1S $T=388740 1001400 0 0 $X=388740 $Y=1001020
X126 2432 2 2427 1 INV1S $T=391220 961080 1 180 $X=389980 $Y=960700
X127 192 2 217 1 INV1S $T=397420 920760 0 0 $X=397420 $Y=920380
X128 2449 2 2484 1 INV1S $T=398040 951000 1 0 $X=398040 $Y=945580
X129 2468 2 2491 1 INV1S $T=398660 971160 0 0 $X=398660 $Y=970780
X130 2497 2 2479 1 INV1S $T=401760 961080 0 180 $X=400520 $Y=955660
X131 2557 2 2562 1 INV1S $T=410440 920760 1 0 $X=410440 $Y=915340
X132 2505 2 2568 1 INV1S $T=411680 930840 0 0 $X=411680 $Y=930460
X133 2542 2 2577 1 INV1S $T=412920 920760 1 0 $X=412920 $Y=915340
X134 2590 2 2578 1 INV1S $T=414780 951000 1 180 $X=413540 $Y=950620
X135 2583 2 2602 1 INV1S $T=414780 951000 1 0 $X=414780 $Y=945580
X136 2593 2 2576 1 INV1S $T=417260 940920 1 180 $X=416020 $Y=940540
X137 2609 2 2616 1 INV1S $T=418500 940920 0 0 $X=418500 $Y=940540
X138 2636 2 2627 1 INV1S $T=421600 940920 0 180 $X=420360 $Y=935500
X139 2640 2 2646 1 INV1S $T=422840 930840 1 0 $X=422840 $Y=925420
X140 2664 2 2655 1 INV1S $T=426560 920760 1 180 $X=425320 $Y=920380
X141 2672 2 2411 1 INV1S $T=428420 1021560 0 180 $X=427180 $Y=1016140
X142 2678 2 2671 1 INV1S $T=429040 920760 1 180 $X=427800 $Y=920380
X143 2672 2 2675 1 INV1S $T=430280 1011480 1 0 $X=430280 $Y=1006060
X144 2744 2 2735 1 INV1S $T=440200 1031640 0 180 $X=438960 $Y=1026220
X145 2735 2 2486 1 INV1S $T=441440 1041720 0 180 $X=440200 $Y=1036300
X146 2735 2 2738 1 INV1S $T=441440 1041720 1 0 $X=441440 $Y=1036300
X147 2750 2 205 1 INV1S $T=442680 1082040 0 180 $X=441440 $Y=1076620
X148 2749 2 227 1 INV1S $T=443300 1041720 1 180 $X=442060 $Y=1041340
X149 2771 2 241 1 INV1S $T=445780 1041720 1 180 $X=444540 $Y=1041340
X150 267 2 2749 1 INV1S $T=445160 1021560 1 0 $X=445160 $Y=1016140
X151 2785 2 2515 1 INV1S $T=448260 1001400 0 180 $X=447020 $Y=995980
X152 2785 2 2549 1 INV1S $T=448260 1001400 1 180 $X=447020 $Y=1001020
X153 2749 2 2790 1 INV1S $T=448260 1061880 0 0 $X=448260 $Y=1061500
X154 2549 2 2799 1 INV1S $T=448880 1011480 1 0 $X=448880 $Y=1006060
X155 2771 2 2800 1 INV1S $T=453220 1051800 0 180 $X=451980 $Y=1046380
X156 2823 2 2672 1 INV1S $T=453840 1001400 1 180 $X=452600 $Y=1001020
X157 2819 2 2771 1 INV1S $T=454460 1051800 0 180 $X=453220 $Y=1046380
X158 280 2 2806 1 INV1S $T=456940 1082040 1 180 $X=455700 $Y=1081660
X159 2860 2 266 1 INV1S $T=459420 920760 0 180 $X=458180 $Y=915340
X160 2750 2 2851 1 INV1S $T=459420 1001400 0 0 $X=459420 $Y=1001020
X161 2867 2 2782 1 INV1S $T=462520 940920 0 180 $X=461280 $Y=935500
X162 290 2 2728 1 INV1S $T=462520 1021560 0 180 $X=461280 $Y=1016140
X163 293 2 294 1 INV1S $T=463760 900600 0 0 $X=463760 $Y=900220
X164 2867 2 2645 1 INV1S $T=464380 1021560 1 0 $X=464380 $Y=1016140
X165 2869 2 2898 1 INV1S $T=468720 1071960 0 0 $X=468720 $Y=1071580
X166 290 2 2908 1 INV1S $T=471820 991320 0 0 $X=471820 $Y=990940
X167 2730 2 2925 1 INV1S $T=473680 940920 0 0 $X=473680 $Y=940540
X168 2926 2 2876 1 INV1S $T=474920 1051800 1 180 $X=473680 $Y=1051420
X169 2806 2 2926 1 INV1S $T=473680 1061880 1 0 $X=473680 $Y=1056460
X170 2926 2 2944 1 INV1S $T=476780 1061880 0 0 $X=476780 $Y=1061500
X171 2961 2 2825 1 INV1S $T=479880 971160 1 180 $X=478640 $Y=970780
X172 2941 2 2961 1 INV1S $T=481740 961080 0 180 $X=480500 $Y=955660
X173 2961 2 2970 1 INV1S $T=480500 971160 0 0 $X=480500 $Y=970780
X174 2971 2 2875 1 INV1S $T=482360 951000 0 180 $X=481120 $Y=945580
X175 2961 2 2955 1 INV1S $T=481120 981240 1 0 $X=481120 $Y=975820
X176 2993 2 2785 1 INV1S $T=485460 1001400 0 180 $X=484220 $Y=995980
X177 2971 2 2941 1 INV1S $T=487320 951000 1 0 $X=487320 $Y=945580
X178 2929 2 3027 1 INV1S $T=491040 1041720 1 0 $X=491040 $Y=1036300
X179 3031 2 2867 1 INV1S $T=492900 940920 0 180 $X=491660 $Y=935500
X180 3026 2 3030 1 INV1S $T=491660 1031640 1 0 $X=491660 $Y=1026220
X181 2807 2 2971 1 INV1S $T=493520 951000 0 180 $X=492280 $Y=945580
X182 2860 2 3060 1 INV1S $T=502200 910680 0 0 $X=502200 $Y=910300
X183 3008 2 3080 1 INV1S $T=502200 1051800 1 0 $X=502200 $Y=1046380
X184 3088 2 3069 1 INV1S $T=504060 971160 0 180 $X=502820 $Y=965740
X185 3095 2 2942 1 INV1S $T=506540 961080 0 180 $X=505300 $Y=955660
X186 3093 2 2993 1 INV1S $T=506540 1001400 1 180 $X=505300 $Y=1001020
X187 3101 2 2860 1 INV1S $T=507160 910680 0 180 $X=505920 $Y=905260
X188 3104 2 3031 1 INV1S $T=507780 940920 0 180 $X=506540 $Y=935500
X189 345 2 2807 1 INV1S $T=508400 920760 1 180 $X=507160 $Y=920380
X190 3122 2 2823 1 INV1S $T=509020 1001400 0 180 $X=507780 $Y=995980
X191 3079 2 345 1 INV1S $T=510880 981240 1 180 $X=509640 $Y=980860
X192 3126 2 3118 1 INV1S $T=511500 1031640 1 180 $X=510260 $Y=1031260
X193 3149 2 3132 1 INV1S $T=515840 961080 1 0 $X=515840 $Y=955660
X194 3149 2 3106 1 INV1S $T=517080 1001400 0 180 $X=515840 $Y=995980
X195 3146 2 3149 1 INV1S $T=517700 951000 1 180 $X=516460 $Y=950620
X196 361 2 3139 1 INV1S $T=522040 910680 1 180 $X=520800 $Y=910300
X197 3213 2 3134 1 INV1S $T=527620 951000 0 180 $X=526380 $Y=945580
X198 3213 2 3228 1 INV1S $T=529480 940920 0 0 $X=529480 $Y=940540
X199 375 2 2990 1 INV1S $T=532580 1031640 1 0 $X=532580 $Y=1026220
X200 3213 2 3258 1 INV1S $T=535060 940920 0 0 $X=535060 $Y=940540
X201 3253 2 3223 1 INV1S $T=536300 981240 0 180 $X=535060 $Y=975820
X202 3255 2 3127 1 INV1S $T=536300 1041720 0 180 $X=535060 $Y=1036300
X203 375 2 383 1 INV1S $T=535680 920760 0 0 $X=535680 $Y=920380
X204 3223 2 3213 1 INV1S $T=535680 951000 0 0 $X=535680 $Y=950620
X205 3255 2 3245 1 INV1S $T=536920 1011480 1 180 $X=535680 $Y=1011100
X206 3301 2 3240 1 INV1S $T=541880 971160 0 180 $X=540640 $Y=965740
X207 3290 2 3255 1 INV1S $T=542500 1011480 0 180 $X=541260 $Y=1006060
X208 395 2 3077 1 INV1S $T=544980 900600 1 180 $X=543740 $Y=900220
X209 3314 2 3146 1 INV1S $T=545600 951000 0 180 $X=544360 $Y=945580
X210 3318 2 3297 1 INV1S $T=546220 910680 0 180 $X=544980 $Y=905260
X211 3334 2 3309 1 INV1S $T=549320 1031640 1 180 $X=548080 $Y=1031260
X212 3334 2 3195 1 INV1S $T=549940 1041720 0 180 $X=548700 $Y=1036300
X213 3348 2 3336 1 INV1S $T=551180 971160 0 0 $X=551180 $Y=970780
X214 3368 2 3334 1 INV1S $T=555520 1031640 1 180 $X=554280 $Y=1031260
X215 3258 2 3372 1 INV1S $T=554900 930840 0 0 $X=554900 $Y=930460
X216 3374 2 3345 1 INV1S $T=556760 1031640 1 180 $X=555520 $Y=1031260
X217 3372 2 3294 1 INV1S $T=558000 930840 1 180 $X=556760 $Y=930460
X218 413 2 3348 1 INV1S $T=559240 971160 1 0 $X=559240 $Y=965740
X219 3372 2 3397 1 INV1S $T=559860 930840 0 0 $X=559860 $Y=930460
X220 3398 2 3303 1 INV1S $T=561100 1001400 0 180 $X=559860 $Y=995980
X221 3400 2 3413 1 INV1S $T=560480 1071960 0 0 $X=560480 $Y=1071580
X222 3343 2 3398 1 INV1S $T=562960 981240 1 180 $X=561720 $Y=980860
X223 3409 2 3374 1 INV1S $T=562960 1041720 0 180 $X=561720 $Y=1036300
X224 3374 2 412 1 INV1S $T=561720 1082040 1 0 $X=561720 $Y=1076620
X225 3413 2 3192 1 INV1S $T=562960 1061880 1 0 $X=562960 $Y=1056460
X226 3348 2 384 1 INV1S $T=564200 971160 0 0 $X=564200 $Y=970780
X227 3311 2 3441 1 INV1S $T=566060 981240 1 0 $X=566060 $Y=975820
X228 3443 2 434 1 INV1S $T=568540 1061880 0 180 $X=567300 $Y=1056460
X229 3398 2 3458 1 INV1S $T=569780 991320 1 0 $X=569780 $Y=985900
X230 3441 2 3377 1 INV1S $T=577840 961080 1 0 $X=577840 $Y=955660
X231 3531 2 3496 1 INV1S $T=586520 971160 1 180 $X=585280 $Y=970780
X232 3535 2 3229 1 INV1S $T=586520 1051800 1 180 $X=585280 $Y=1051420
X233 3441 2 3532 1 INV1S $T=585900 961080 0 0 $X=585900 $Y=960700
X234 383 2 3535 1 INV1S $T=591480 900600 0 0 $X=591480 $Y=900220
X235 3584 2 3290 1 INV1S $T=598300 940920 1 180 $X=597060 $Y=940540
X236 3606 2 3586 1 INV1S $T=603880 951000 0 180 $X=602640 $Y=945580
X237 496 2 3616 1 INV1S $T=603260 1061880 1 0 $X=603260 $Y=1056460
X238 3535 2 3620 1 INV1S $T=603880 1051800 0 0 $X=603880 $Y=1051420
X239 3623 2 3328 1 INV1S $T=606360 951000 0 180 $X=605120 $Y=945580
X240 3420 2 3628 1 INV1S $T=605740 961080 0 0 $X=605740 $Y=960700
X241 3636 2 3305 1 INV1S $T=607600 961080 0 180 $X=606360 $Y=955660
X242 3602 2 3633 1 INV1S $T=606360 1082040 1 0 $X=606360 $Y=1076620
X243 3401 2 3652 1 INV1S $T=610700 1041720 1 0 $X=610700 $Y=1036300
X244 3652 2 3548 1 INV1S $T=611940 1061880 0 180 $X=610700 $Y=1056460
X245 3685 2 3654 1 INV1S $T=617520 971160 1 180 $X=616280 $Y=970780
X246 3646 2 3582 1 INV1S $T=616280 1021560 0 0 $X=616280 $Y=1021180
X247 3689 2 3666 1 INV1S $T=618140 1082040 0 180 $X=616900 $Y=1076620
X248 3652 2 3697 1 INV1S $T=618760 1041720 0 0 $X=618760 $Y=1041340
X249 3646 2 3730 1 INV1S $T=622480 1021560 0 0 $X=622480 $Y=1021180
X250 3739 2 3752 1 INV1S $T=624960 940920 0 0 $X=624960 $Y=940540
X251 534 2 3765 1 INV1S $T=629300 951000 0 0 $X=629300 $Y=950620
X252 3711 2 3710 1 INV1S $T=631160 991320 1 180 $X=629920 $Y=990940
X253 3628 2 3786 1 INV1S $T=631780 961080 0 0 $X=631780 $Y=960700
X254 3711 2 3753 1 INV1S $T=633640 1011480 1 0 $X=633640 $Y=1006060
X255 3628 2 3834 1 INV1S $T=643560 961080 1 0 $X=643560 $Y=955660
X256 3838 2 3746 1 INV1S $T=645420 1001400 0 180 $X=644180 $Y=995980
X257 3839 2 3838 1 INV1S $T=646040 1001400 1 0 $X=646040 $Y=995980
X258 3838 2 3677 1 INV1S $T=647900 1021560 1 0 $X=647900 $Y=1016140
X259 565 2 3863 1 INV1S $T=649140 1061880 1 0 $X=649140 $Y=1056460
X260 565 2 567 1 INV1S $T=649140 1082040 0 0 $X=649140 $Y=1081660
X261 3865 2 3872 1 INV1S $T=651620 920760 0 0 $X=651620 $Y=920380
X262 3820 2 3878 1 INV1S $T=652240 1082040 1 0 $X=652240 $Y=1076620
X263 577 2 3824 1 INV1S $T=654100 910680 0 180 $X=652860 $Y=905260
X264 3896 2 3795 1 INV1S $T=656580 961080 0 180 $X=655340 $Y=955660
X265 580 2 574 1 INV1S $T=657820 920760 1 180 $X=656580 $Y=920380
X266 3900 2 3629 1 INV1S $T=657820 961080 0 180 $X=656580 $Y=955660
X267 3914 2 3813 1 INV1S $T=659680 1011480 0 180 $X=658440 $Y=1006060
X268 588 2 3903 1 INV1S $T=660920 930840 0 180 $X=659680 $Y=925420
X269 593 2 577 1 INV1S $T=662780 910680 0 180 $X=661540 $Y=905260
X270 585 2 534 1 INV1S $T=661540 940920 1 0 $X=661540 $Y=935500
X271 3947 2 3941 1 INV1S $T=665260 1031640 1 180 $X=664020 $Y=1031260
X272 534 2 3961 1 INV1S $T=665880 951000 1 0 $X=665880 $Y=945580
X273 3951 2 3940 1 INV1S $T=667120 961080 0 180 $X=665880 $Y=955660
X274 3971 2 3867 1 INV1S $T=668360 981240 1 180 $X=667120 $Y=980860
X275 3801 2 3975 1 INV1S $T=667740 951000 1 0 $X=667740 $Y=945580
X276 3980 2 3860 1 INV1S $T=669600 1011480 0 180 $X=668360 $Y=1006060
X277 602 2 3965 1 INV1S $T=669600 1082040 0 180 $X=668360 $Y=1076620
X278 3983 2 3812 1 INV1S $T=670220 951000 0 180 $X=668980 $Y=945580
X279 3984 2 3839 1 INV1S $T=670220 981240 1 180 $X=668980 $Y=980860
X280 580 2 3999 1 INV1S $T=670840 951000 1 0 $X=670840 $Y=945580
X281 3636 2 3962 1 INV1S $T=671460 961080 1 0 $X=671460 $Y=955660
X282 4014 2 3858 1 INV1S $T=673940 1001400 0 180 $X=672700 $Y=995980
X283 610 2 4010 1 INV1S $T=673320 1082040 0 0 $X=673320 $Y=1081660
X284 607 2 3685 1 INV1S $T=677040 951000 0 180 $X=675800 $Y=945580
X285 608 2 3636 1 INV1S $T=677040 951000 1 180 $X=675800 $Y=950620
X286 3685 2 4033 1 INV1S $T=677040 961080 0 0 $X=677040 $Y=960700
X287 4034 2 3852 1 INV1S $T=678280 1082040 0 180 $X=677040 $Y=1076620
X288 620 2 3900 1 INV1S $T=677660 951000 1 0 $X=677660 $Y=945580
X289 621 2 3972 1 INV1S $T=678900 1031640 0 180 $X=677660 $Y=1026220
X290 3316 2 4024 1 INV1S $T=678280 1001400 1 0 $X=678280 $Y=995980
X291 4041 2 582 1 INV1S $T=679520 1082040 0 180 $X=678280 $Y=1076620
X292 3969 2 4034 1 INV1S $T=681380 1082040 0 180 $X=680140 $Y=1076620
X293 3900 2 4054 1 INV1S $T=680760 961080 0 0 $X=680760 $Y=960700
X294 629 2 601 1 INV1S $T=682620 920760 1 180 $X=681380 $Y=920380
X295 4041 2 630 1 INV1S $T=681380 1071960 0 0 $X=681380 $Y=1071580
X296 557 2 4075 1 INV1S $T=682000 930840 1 0 $X=682000 $Y=925420
X297 626 2 4069 1 INV1S $T=683240 920760 0 0 $X=683240 $Y=920380
X298 4069 2 3891 1 INV1S $T=686340 961080 0 180 $X=685100 $Y=955660
X299 4116 2 4029 1 INV1S $T=691300 991320 1 0 $X=691300 $Y=985900
X300 4125 2 4113 1 INV1S $T=693160 1071960 1 180 $X=691920 $Y=1071580
X301 4069 2 4126 1 INV1S $T=692540 961080 1 0 $X=692540 $Y=955660
X302 4024 2 4128 1 INV1S $T=692540 1001400 0 0 $X=692540 $Y=1001020
X303 4034 2 4131 1 INV1S $T=693160 1071960 0 0 $X=693160 $Y=1071580
X304 3971 2 4137 1 INV1S $T=695020 1001400 0 0 $X=695020 $Y=1001020
X305 4146 2 3971 1 INV1S $T=697500 991320 0 180 $X=696260 $Y=985900
X306 4150 2 3832 1 INV1S $T=698120 1051800 1 180 $X=696880 $Y=1051420
X307 4142 2 650 1 INV1S $T=696880 1082040 0 0 $X=696880 $Y=1081660
X308 4154 2 4159 1 INV1S $T=698120 1041720 1 0 $X=698120 $Y=1036300
X309 4158 2 4150 1 INV1S $T=699360 1051800 0 180 $X=698120 $Y=1046380
X310 4019 2 4142 1 INV1S $T=698740 1071960 0 0 $X=698740 $Y=1071580
X311 4029 2 4154 1 INV1S $T=701220 1031640 1 180 $X=699980 $Y=1031260
X312 4075 2 4180 1 INV1S $T=701220 930840 1 0 $X=701220 $Y=925420
X313 638 2 4184 1 INV1S $T=701220 1082040 0 0 $X=701220 $Y=1081660
X314 4103 2 656 1 INV1S $T=704320 1071960 1 180 $X=703080 $Y=1071580
X315 659 2 3096 1 INV1S $T=704940 951000 0 180 $X=703700 $Y=945580
X316 4128 2 4064 1 INV1S $T=706180 1001400 0 180 $X=704940 $Y=995980
X317 4219 2 4055 1 INV1S $T=709280 1011480 1 180 $X=708040 $Y=1011100
X318 4142 2 4221 1 INV1S $T=709280 1071960 0 0 $X=709280 $Y=1071580
X319 4128 2 4217 1 INV1S $T=709900 1001400 1 0 $X=709900 $Y=995980
X320 3747 2 4240 1 INV1S $T=711760 1011480 0 0 $X=711760 $Y=1011100
X321 4241 2 3947 1 INV1S $T=713000 1031640 1 180 $X=711760 $Y=1031260
X322 4246 2 651 1 INV1S $T=714240 910680 0 180 $X=713000 $Y=905260
X323 4153 2 4246 1 INV1S $T=713000 920760 1 0 $X=713000 $Y=915340
X324 4226 2 4241 1 INV1S $T=713620 991320 1 0 $X=713620 $Y=985900
X325 4191 2 4236 1 INV1S $T=713620 1021560 1 0 $X=713620 $Y=1016140
X326 4246 2 4232 1 INV1S $T=714240 910680 1 0 $X=714240 $Y=905260
X327 4219 2 4149 1 INV1S $T=716720 1021560 1 0 $X=716720 $Y=1016140
X328 669 2 4260 1 INV1S $T=716720 1082040 0 0 $X=716720 $Y=1081660
X329 4263 2 3623 1 INV1S $T=719200 951000 0 180 $X=717960 $Y=945580
X330 4241 2 4271 1 INV1S $T=719200 1031640 0 0 $X=719200 $Y=1031260
X331 4191 2 4273 1 INV1S $T=719820 1021560 1 0 $X=719820 $Y=1016140
X332 4281 2 4087 1 INV1S $T=722300 951000 1 180 $X=721060 $Y=950620
X333 4116 2 4278 1 INV1S $T=721680 1031640 1 0 $X=721680 $Y=1026220
X334 3623 2 4288 1 INV1S $T=722300 951000 0 0 $X=722300 $Y=950620
X335 4300 2 4141 1 INV1S $T=723540 1011480 0 180 $X=722300 $Y=1006060
X336 4240 2 667 1 INV1S $T=724160 1011480 1 180 $X=722920 $Y=1011100
X337 4297 2 4219 1 INV1S $T=724780 981240 0 180 $X=723540 $Y=975820
X338 4306 2 4291 1 INV1S $T=726020 991320 1 180 $X=724780 $Y=990940
X339 4307 2 4300 1 INV1S $T=726020 1011480 0 180 $X=724780 $Y=1006060
X340 483 2 688 1 INV1S $T=725400 910680 1 0 $X=725400 $Y=905260
X341 4253 2 4313 1 INV1S $T=725400 991320 1 0 $X=725400 $Y=985900
X342 4300 2 4308 1 INV1S $T=726020 1011480 0 0 $X=726020 $Y=1011100
X343 659 2 4324 1 INV1S $T=726640 951000 1 0 $X=726640 $Y=945580
X344 529 2 4331 1 INV1S $T=728500 951000 1 0 $X=728500 $Y=945580
X345 4331 2 4340 1 INV1S $T=728500 951000 0 0 $X=728500 $Y=950620
X346 4306 2 4230 1 INV1S $T=730980 1011480 0 0 $X=730980 $Y=1011100
X347 4366 2 4171 1 INV1S $T=733460 1001400 0 180 $X=732220 $Y=995980
X348 4364 2 4338 1 INV1S $T=733460 1082040 0 180 $X=732220 $Y=1076620
X349 4322 2 4297 1 INV1S $T=732840 971160 1 0 $X=732840 $Y=965740
X350 4331 2 4368 1 INV1S $T=733460 951000 1 0 $X=733460 $Y=945580
X351 4353 2 4366 1 INV1S $T=733460 991320 0 0 $X=733460 $Y=990940
X352 4366 2 4357 1 INV1S $T=733460 1001400 1 0 $X=733460 $Y=995980
X353 4381 2 4306 1 INV1S $T=736560 991320 0 180 $X=735320 $Y=985900
X354 700 2 4365 1 INV1S $T=736560 920760 0 0 $X=736560 $Y=920380
X355 4387 2 4378 1 INV1S $T=737800 981240 0 180 $X=736560 $Y=975820
X356 705 2 4387 1 INV1S $T=737800 981240 1 0 $X=737800 $Y=975820
X357 4313 2 4408 1 INV1S $T=740900 991320 1 0 $X=740900 $Y=985900
X358 4313 2 4332 1 INV1S $T=741520 981240 0 0 $X=741520 $Y=980860
X359 710 2 3086 1 INV1S $T=743380 951000 1 0 $X=743380 $Y=945580
X360 4418 2 4307 1 INV1S $T=745240 991320 0 180 $X=744000 $Y=985900
X361 4240 2 4432 1 INV1S $T=747100 1011480 0 0 $X=747100 $Y=1011100
X362 4421 2 4442 1 INV1S $T=748340 1021560 1 0 $X=748340 $Y=1016140
X363 3316 2 4459 1 INV1S $T=752060 991320 0 0 $X=752060 $Y=990940
X364 4268 2 4473 1 INV1S $T=752680 1071960 0 0 $X=752680 $Y=1071580
X365 4459 2 4490 1 INV1S $T=757640 991320 1 0 $X=757640 $Y=985900
X366 726 2 4441 1 INV1S $T=758260 951000 0 0 $X=758260 $Y=950620
X367 4473 2 731 1 INV1S $T=764460 1082040 1 0 $X=764460 $Y=1076620
X368 4490 2 4466 1 INV1S $T=766320 971160 0 180 $X=765080 $Y=965740
X369 739 2 717 1 INV1S $T=766320 900600 0 0 $X=766320 $Y=900220
X370 4442 2 4531 1 INV1S $T=768180 1021560 1 0 $X=768180 $Y=1016140
X371 4546 2 4528 1 INV1S $T=769420 1031640 0 180 $X=768180 $Y=1026220
X372 4075 2 4545 1 INV1S $T=770040 910680 0 180 $X=768800 $Y=905260
X373 4532 2 4546 1 INV1S $T=770660 1031640 0 180 $X=769420 $Y=1026220
X374 4546 2 4522 1 INV1S $T=769420 1041720 0 0 $X=769420 $Y=1041340
X375 4442 2 4562 1 INV1S $T=770040 1021560 1 0 $X=770040 $Y=1016140
X376 711 2 4571 1 INV1S $T=771280 1071960 0 0 $X=771280 $Y=1071580
X377 4544 2 4575 1 INV1S $T=771900 1071960 1 0 $X=771900 $Y=1066540
X378 758 2 4607 1 INV1S $T=775000 900600 0 0 $X=775000 $Y=900220
X379 4601 2 4593 1 INV1S $T=776860 1001400 1 180 $X=775620 $Y=1001020
X380 4490 2 4621 1 INV1S $T=778720 971160 0 0 $X=778720 $Y=970780
X381 4490 2 4478 1 INV1S $T=779340 991320 1 0 $X=779340 $Y=985900
X382 4627 2 4511 1 INV1S $T=780580 1041720 1 180 $X=779340 $Y=1041340
X383 4604 2 4627 1 INV1S $T=779340 1061880 0 0 $X=779340 $Y=1061500
X384 4607 2 4633 1 INV1S $T=784300 900600 0 0 $X=784300 $Y=900220
X385 4571 2 4673 1 INV1S $T=788020 1071960 0 0 $X=788020 $Y=1071580
X386 4075 2 4717 1 INV1S $T=791120 910680 1 0 $X=791120 $Y=905260
X387 4762 2 4692 1 INV1S $T=799800 961080 0 180 $X=798560 $Y=955660
X388 4621 2 4762 1 INV1S $T=801040 961080 1 180 $X=799800 $Y=960700
X389 4627 2 4766 1 INV1S $T=799800 1061880 1 0 $X=799800 $Y=1056460
X390 4762 2 4781 1 INV1S $T=801040 961080 0 0 $X=801040 $Y=960700
X391 4792 2 4775 1 INV1S $T=804760 1011480 1 0 $X=804760 $Y=1006060
X392 4806 2 4794 1 INV1S $T=806620 940920 0 180 $X=805380 $Y=935500
X393 4822 2 4829 1 INV1S $T=807860 1041720 0 0 $X=807860 $Y=1041340
X394 785 2 4830 1 INV1S $T=808480 910680 0 0 $X=808480 $Y=910300
X395 4793 2 4809 1 INV1S $T=808480 1021560 1 0 $X=808480 $Y=1016140
X396 4806 2 4780 1 INV1S $T=809720 940920 1 0 $X=809720 $Y=935500
X397 779 2 4797 1 INV1S $T=812200 1021560 0 180 $X=810960 $Y=1016140
X398 4800 2 4832 1 INV1S $T=812200 1061880 0 180 $X=810960 $Y=1056460
X399 4695 2 4806 1 INV1S $T=812820 940920 1 180 $X=811580 $Y=940540
X400 4850 2 4795 1 INV1S $T=812820 981240 0 180 $X=811580 $Y=975820
X401 4751 2 4837 1 INV1S $T=811580 1011480 1 0 $X=811580 $Y=1006060
X402 4850 2 4803 1 INV1S $T=812200 971160 1 0 $X=812200 $Y=965740
X403 836 2 4861 1 INV1S $T=815920 910680 0 180 $X=814680 $Y=905260
X404 4830 2 4871 1 INV1S $T=814680 920760 0 0 $X=814680 $Y=920380
X405 4852 2 4872 1 INV1S $T=814680 1011480 0 0 $X=814680 $Y=1011100
X406 4781 2 4888 1 INV1S $T=817780 961080 0 0 $X=817780 $Y=960700
X407 4890 2 4853 1 INV1S $T=819020 1001400 0 180 $X=817780 $Y=995980
X408 4902 2 4850 1 INV1S $T=821500 961080 0 180 $X=820260 $Y=955660
X409 4879 2 4897 1 INV1S $T=822120 910680 1 180 $X=820880 $Y=910300
X410 4888 2 4908 1 INV1S $T=822740 961080 1 0 $X=822740 $Y=955660
X411 4888 2 4909 1 INV1S $T=824600 971160 1 0 $X=824600 $Y=965740
X412 853 2 4600 1 INV1S $T=827080 930840 0 0 $X=827080 $Y=930460
X413 4927 2 4902 1 INV1S $T=828320 961080 0 180 $X=827080 $Y=955660
X414 4856 2 4931 1 INV1S $T=827080 1021560 1 0 $X=827080 $Y=1016140
X415 4931 2 4778 1 INV1S $T=828940 1001400 0 180 $X=827700 $Y=995980
X416 4931 2 4935 1 INV1S $T=828940 1011480 1 0 $X=828940 $Y=1006060
X417 4931 2 4942 1 INV1S $T=828940 1011480 0 0 $X=828940 $Y=1011100
X418 4473 2 4951 1 INV1S $T=832660 1082040 0 180 $X=831420 $Y=1076620
X419 4473 2 861 1 INV1S $T=832660 1082040 1 0 $X=832660 $Y=1076620
X420 4926 2 4967 1 INV1S $T=833900 951000 0 0 $X=833900 $Y=950620
X421 5004 2 4611 1 INV1S $T=841960 971160 0 180 $X=840720 $Y=965740
X422 5004 2 5009 1 INV1S $T=841340 981240 1 0 $X=841340 $Y=975820
X423 5006 2 4952 1 INV1S $T=842580 991320 1 180 $X=841340 $Y=990940
X424 4990 2 5007 1 INV1S $T=841340 1011480 0 0 $X=841340 $Y=1011100
X425 872 2 5004 1 INV1S $T=843200 951000 0 180 $X=841960 $Y=945580
X426 5027 2 5000 1 INV1S $T=845680 981240 1 180 $X=844440 $Y=980860
X427 4951 2 5042 1 INV1S $T=845060 1041720 0 0 $X=845060 $Y=1041340
X428 4924 2 5037 1 INV1S $T=845680 991320 1 0 $X=845680 $Y=985900
X429 4883 2 5046 1 INV1S $T=846920 1031640 1 0 $X=846920 $Y=1026220
X430 5042 2 5031 1 INV1S $T=846920 1041720 0 0 $X=846920 $Y=1041340
X431 5037 2 5050 1 INV1S $T=847540 991320 1 0 $X=847540 $Y=985900
X432 5042 2 5064 1 INV1S $T=849400 1041720 0 0 $X=849400 $Y=1041340
X433 4607 2 4606 1 INV1S $T=855600 1021560 0 0 $X=855600 $Y=1021180
X434 5000 2 5099 1 INV1S $T=856220 991320 1 0 $X=856220 $Y=985900
X435 5098 2 5108 1 INV1S $T=857460 940920 0 0 $X=857460 $Y=940540
X436 862 2 899 1 INV1S $T=863040 1082040 0 0 $X=863040 $Y=1081660
X437 5070 2 5162 1 INV1S $T=866140 930840 0 0 $X=866140 $Y=930460
X438 5162 2 906 1 INV1S $T=869240 940920 1 0 $X=869240 $Y=935500
X439 5155 2 5177 1 INV1S $T=869240 1041720 1 0 $X=869240 $Y=1036300
X440 5183 2 5132 1 INV1S $T=871720 1031640 1 180 $X=870480 $Y=1031260
X441 5182 2 5196 1 INV1S $T=871100 981240 1 0 $X=871100 $Y=975820
X442 5031 2 5183 1 INV1S $T=871720 1031640 0 0 $X=871720 $Y=1031260
X443 4134 2 5182 1 INV1S $T=872960 1001400 1 0 $X=872960 $Y=995980
X444 5041 2 5213 1 INV1S $T=874200 1021560 0 0 $X=874200 $Y=1021180
X445 5099 2 5224 1 INV1S $T=876060 981240 0 0 $X=876060 $Y=980860
X446 4571 2 918 1 INV1S $T=881640 1082040 1 180 $X=880400 $Y=1081660
X447 4571 2 924 1 INV1S $T=881640 1082040 0 0 $X=881640 $Y=1081660
X448 5099 2 5263 1 INV1S $T=882260 981240 0 0 $X=882260 $Y=980860
X449 5269 2 5274 1 INV1S $T=884120 1011480 1 0 $X=884120 $Y=1006060
X450 5274 2 5275 1 INV1S $T=884740 1021560 0 0 $X=884740 $Y=1021180
X451 5280 2 5200 1 INV1S $T=886600 940920 0 180 $X=885360 $Y=935500
X452 5249 2 5296 1 INV1S $T=885980 1011480 1 0 $X=885980 $Y=1006060
X453 5274 2 5245 1 INV1S $T=885980 1031640 0 0 $X=885980 $Y=1031260
X454 5327 2 5318 1 INV1S $T=893420 1011480 0 180 $X=892180 $Y=1006060
X455 5287 2 5280 1 INV1S $T=892800 951000 1 0 $X=892800 $Y=945580
X456 5296 2 5331 1 INV1S $T=892800 1011480 0 0 $X=892800 $Y=1011100
X457 5331 2 5149 1 INV1S $T=894660 1041720 0 180 $X=893420 $Y=1036300
X458 5331 2 5353 1 INV1S $T=897140 1011480 1 0 $X=897140 $Y=1006060
X459 945 2 938 1 INV1S $T=898380 1082040 0 0 $X=898380 $Y=1081660
X460 5367 2 5359 1 INV1S $T=900240 1011480 1 180 $X=899000 $Y=1011100
X461 5255 2 5435 1 INV1S $T=912020 940920 0 0 $X=912020 $Y=940540
X462 5340 2 5420 1 INV1S $T=912020 981240 0 0 $X=912020 $Y=980860
X463 5420 2 5432 1 INV1S $T=923180 991320 1 180 $X=921940 $Y=990940
X464 5420 2 5451 1 INV1S $T=925040 991320 1 180 $X=923800 $Y=990940
X465 5485 2 5490 1 INV1S $T=925660 951000 1 0 $X=925660 $Y=945580
X466 5420 2 5487 1 INV1S $T=926900 991320 1 0 $X=926900 $Y=985900
X467 999 2 5505 1 INV1S $T=928760 920760 0 0 $X=928760 $Y=920380
X468 5420 2 5503 1 INV1S $T=928760 991320 1 0 $X=928760 $Y=985900
X469 5505 2 5508 1 INV1S $T=930620 971160 0 0 $X=930620 $Y=970780
X470 5535 2 5537 1 INV1S $T=933720 951000 1 0 $X=933720 $Y=945580
X471 688 2 5576 1 INV1S $T=937440 920760 1 0 $X=937440 $Y=915340
X472 1011 2 5553 1 INV1S $T=937440 940920 1 0 $X=937440 $Y=935500
X473 5499 2 5603 1 INV1S $T=939920 951000 0 0 $X=939920 $Y=950620
X474 1011 2 5545 1 INV1S $T=941160 1011480 0 180 $X=939920 $Y=1006060
X475 5571 2 1021 1 INV1S $T=940540 930840 0 0 $X=940540 $Y=930460
X476 5533 2 5610 1 INV1S $T=945500 951000 0 0 $X=945500 $Y=950620
X477 5526 2 5656 1 INV1S $T=951080 991320 0 0 $X=951080 $Y=990940
X478 5683 2 5575 1 INV1S $T=957280 1071960 0 180 $X=956040 $Y=1066540
X479 5663 2 5669 1 INV1S $T=956660 940920 0 0 $X=956660 $Y=940540
X480 5433 2 5764 1 INV1S $T=970920 1061880 0 0 $X=970920 $Y=1061500
X481 5764 2 5746 1 INV1S $T=975880 1061880 1 180 $X=974640 $Y=1061500
X482 5182 2 5717 1 INV1S $T=979600 1011480 1 180 $X=978360 $Y=1011100
X483 5182 2 5790 1 INV1S $T=983320 961080 1 0 $X=983320 $Y=955660
X484 5853 2 5858 1 INV1S $T=993240 971160 0 0 $X=993240 $Y=970780
X485 5790 2 5860 1 INV1S $T=993860 930840 1 0 $X=993860 $Y=925420
X486 5856 2 5853 1 INV1S $T=993860 961080 1 0 $X=993860 $Y=955660
X487 5853 2 5857 1 INV1S $T=995100 991320 1 180 $X=993860 $Y=990940
X488 5860 2 5682 1 INV1S $T=996960 930840 0 180 $X=995720 $Y=925420
X489 5860 2 5765 1 INV1S $T=998820 930840 1 0 $X=998820 $Y=925420
X490 1100 2 5887 1 INV1S $T=1003780 1001400 1 180 $X=1002540 $Y=1001020
X491 5907 2 5905 1 INV1S $T=1003780 940920 1 0 $X=1003780 $Y=935500
X492 5911 2 5918 1 INV1S $T=1003780 981240 1 0 $X=1003780 $Y=975820
X493 5911 2 5897 1 INV1S $T=1005640 991320 0 180 $X=1004400 $Y=985900
X494 5930 2 5911 1 INV1S $T=1006260 961080 0 180 $X=1005020 $Y=955660
X495 5860 2 5938 1 INV1S $T=1006260 930840 0 0 $X=1006260 $Y=930460
X496 5958 2 1109 1 INV1S $T=1009980 940920 0 180 $X=1008740 $Y=935500
X497 5486 2 5958 1 INV1S $T=1012460 940920 1 180 $X=1011220 $Y=940540
X498 1126 2 5921 1 INV1S $T=1013700 910680 1 0 $X=1013700 $Y=905260
X499 1134 2 6002 1 INV1S $T=1018040 1011480 1 0 $X=1018040 $Y=1006060
X500 5922 2 6020 1 INV1S $T=1019280 1021560 1 0 $X=1019280 $Y=1016140
X501 6014 2 6024 1 INV1S $T=1021760 1001400 1 0 $X=1021760 $Y=995980
X502 6031 2 1135 1 INV1S $T=1023620 1071960 0 180 $X=1022380 $Y=1066540
X503 5497 2 6046 1 INV1S $T=1026720 991320 0 0 $X=1026720 $Y=990940
X504 6050 2 6045 1 INV1S $T=1028580 940920 1 180 $X=1027340 $Y=940540
X505 6076 2 6078 1 INV1S $T=1032300 971160 1 0 $X=1032300 $Y=965740
X506 6075 2 6081 1 INV1S $T=1032920 951000 1 0 $X=1032920 $Y=945580
X507 6045 2 6082 1 INV1S $T=1032920 971160 0 0 $X=1032920 $Y=970780
X508 6082 2 6063 1 INV1S $T=1035400 981240 1 180 $X=1034160 $Y=980860
X509 6082 2 6080 1 INV1S $T=1035400 991320 1 0 $X=1035400 $Y=985900
X510 6018 2 6105 1 INV1S $T=1036640 910680 0 0 $X=1036640 $Y=910300
X511 6105 2 1161 1 INV1S $T=1037260 920760 1 0 $X=1037260 $Y=915340
X512 6039 2 6111 1 INV1S $T=1037880 951000 0 0 $X=1037880 $Y=950620
X513 6046 2 5983 1 INV1S $T=1037880 1001400 0 0 $X=1037880 $Y=1001020
X514 5182 2 6093 1 INV1S $T=1038500 1031640 1 0 $X=1038500 $Y=1026220
X515 6111 2 6101 1 INV1S $T=1039740 971160 1 0 $X=1039740 $Y=965740
X516 6150 2 6158 1 INV1S $T=1045940 1011480 0 0 $X=1045940 $Y=1011100
X517 6150 2 1169 1 INV1S $T=1048420 1031640 1 180 $X=1047180 $Y=1031260
X518 6142 2 6150 1 INV1S $T=1049040 1011480 0 180 $X=1047800 $Y=1006060
X519 1180 2 6141 1 INV1S $T=1049040 951000 1 0 $X=1049040 $Y=945580
X520 6185 2 6181 1 INV1S $T=1054620 951000 0 0 $X=1054620 $Y=950620
X521 6196 2 6190 1 INV1S $T=1057100 951000 1 180 $X=1055860 $Y=950620
X522 1126 2 1193 1 INV1S $T=1056480 900600 0 0 $X=1056480 $Y=900220
X523 6211 2 6231 1 INV1S $T=1061440 951000 1 0 $X=1061440 $Y=945580
X524 1180 2 6223 1 INV1S $T=1061440 951000 0 0 $X=1061440 $Y=950620
X525 6230 2 1198 1 INV1S $T=1065160 1041720 0 180 $X=1063920 $Y=1036300
X526 6249 2 6241 1 INV1S $T=1065780 1001400 0 180 $X=1064540 $Y=995980
X527 6300 2 6146 1 INV1S $T=1076320 940920 0 180 $X=1075080 $Y=935500
X528 1216 2 6304 1 INV1S $T=1076940 1011480 0 0 $X=1076940 $Y=1011100
X529 6167 2 6300 1 INV1S $T=1078800 930840 0 180 $X=1077560 $Y=925420
X530 6300 2 6162 1 INV1S $T=1077560 940920 0 0 $X=1077560 $Y=940540
X531 6261 2 1214 1 INV1S $T=1080040 910680 0 0 $X=1080040 $Y=910300
X532 6046 2 6316 1 INV1S $T=1086240 1001400 0 180 $X=1085000 $Y=995980
X533 6354 2 6336 1 INV1S $T=1088720 951000 1 180 $X=1087480 $Y=950620
X534 6312 2 6354 1 INV1S $T=1088100 940920 0 0 $X=1088100 $Y=940540
X535 6046 2 6399 1 INV1S $T=1100500 1001400 0 180 $X=1099260 $Y=995980
X536 6046 2 6468 1 INV1S $T=1109800 991320 1 0 $X=1109800 $Y=985900
X537 1247 2 6488 1 INV1S $T=1112280 991320 1 0 $X=1112280 $Y=985900
X538 1274 2 1286 1 INV1S $T=1126540 930840 0 0 $X=1126540 $Y=930460
X539 1286 2 1287 1 INV1S $T=1128400 900600 0 0 $X=1128400 $Y=900220
X540 1286 2 6532 1 INV1S $T=1128400 1001400 0 0 $X=1128400 $Y=1001020
X541 5 1 2 3 BUF1S $T=223200 930840 1 180 $X=220720 $Y=930460
X542 1388 1 2 1326 BUF1S $T=231880 1001400 0 180 $X=229400 $Y=995980
X543 1402 1 2 1417 BUF1S $T=234980 1011480 0 0 $X=234980 $Y=1011100
X544 1451 1 2 1358 BUF1S $T=243040 1001400 0 180 $X=240560 $Y=995980
X545 1509 1 2 1388 BUF1S $T=251100 1001400 0 180 $X=248620 $Y=995980
X546 27 1 2 1576 BUF1S $T=258540 940920 1 0 $X=258540 $Y=935500
X547 1615 1 2 31 BUF1S $T=266600 940920 1 180 $X=264120 $Y=940540
X548 1618 1 2 1400 BUF1S $T=267220 1001400 0 180 $X=264740 $Y=995980
X549 1608 1 2 1586 BUF1S $T=265360 1011480 0 0 $X=265360 $Y=1011100
X550 1630 1 2 1544 BUF1S $T=269080 1021560 1 180 $X=266600 $Y=1021180
X551 1674 1 2 1378 BUF1S $T=274660 1031640 0 180 $X=272180 $Y=1026220
X552 1554 1 2 1609 BUF1S $T=274040 1011480 0 0 $X=274040 $Y=1011100
X553 1716 1 2 1451 BUF1S $T=280240 1011480 1 180 $X=277760 $Y=1011100
X554 54 1 2 1695 BUF1S $T=278380 940920 1 0 $X=278380 $Y=935500
X555 1754 1 2 1333 BUF1S $T=283340 1031640 1 180 $X=280860 $Y=1031260
X556 1644 1 2 1717 BUF1S $T=280860 1041720 1 0 $X=280860 $Y=1036300
X557 38 1 2 1734 BUF1S $T=282720 940920 1 0 $X=282720 $Y=935500
X558 1689 1 2 1389 BUF1S $T=284580 1041720 1 0 $X=284580 $Y=1036300
X559 1749 1 2 1452 BUF1S $T=287060 1041720 1 180 $X=284580 $Y=1041340
X560 1800 1 2 1403 BUF1S $T=288920 1031640 0 180 $X=286440 $Y=1026220
X561 64 1 2 1746 BUF1S $T=292640 920760 0 180 $X=290160 $Y=915340
X562 1799 1 2 1509 BUF1S $T=292640 1001400 0 180 $X=290160 $Y=995980
X563 1609 1 2 1808 BUF1S $T=292020 1041720 0 0 $X=292020 $Y=1041340
X564 1796 1 2 1807 BUF1S $T=292640 1001400 0 0 $X=292640 $Y=1001020
X565 72 1 2 76 BUF1S $T=298840 991320 0 0 $X=298840 $Y=990940
X566 77 1 2 1772 BUF1S $T=303180 951000 1 180 $X=300700 $Y=950620
X567 1796 1 2 1800 BUF1S $T=304420 1031640 1 0 $X=304420 $Y=1026220
X568 1912 1 2 1674 BUF1S $T=310000 1031640 0 180 $X=307520 $Y=1026220
X569 93 1 2 1871 BUF1S $T=310000 920760 0 0 $X=310000 $Y=920380
X570 1541 1 2 1913 BUF1S $T=311240 1031640 1 0 $X=311240 $Y=1026220
X571 1939 1 2 1897 BUF1S $T=314340 1001400 1 180 $X=311860 $Y=1001020
X572 106 1 2 1902 BUF1S $T=315580 920760 1 180 $X=313100 $Y=920380
X573 112 1 2 1943 BUF1S $T=318680 940920 0 180 $X=316200 $Y=935500
X574 107 1 2 1906 BUF1S $T=316820 930840 1 0 $X=316820 $Y=925420
X575 108 1 2 1923 BUF1S $T=316820 1021560 1 0 $X=316820 $Y=1016140
X576 1911 1 2 1921 BUF1S $T=318060 930840 0 0 $X=318060 $Y=930460
X577 1880 1 2 1972 BUF1S $T=318060 961080 1 0 $X=318060 $Y=955660
X578 1974 1 2 1778 BUF1S $T=321160 940920 1 180 $X=318680 $Y=940540
X579 75 1 2 1976 BUF1S $T=319300 1021560 1 0 $X=319300 $Y=1016140
X580 1911 1 2 118 BUF1S $T=319920 910680 1 0 $X=319920 $Y=905260
X581 119 1 2 1754 BUF1S $T=322400 1041720 0 180 $X=319920 $Y=1036300
X582 80 1 2 1917 BUF1S $T=320540 920760 0 0 $X=320540 $Y=920380
X583 1968 1 2 110 BUF1S $T=321160 910680 0 0 $X=321160 $Y=910300
X584 1550 1 2 122 BUF1S $T=323640 910680 1 0 $X=323640 $Y=905260
X585 129 1 2 1689 BUF1S $T=329840 1051800 0 180 $X=327360 $Y=1046380
X586 127 1 2 2055 BUF1S $T=328600 910680 1 0 $X=328600 $Y=905260
X587 128 1 2 1874 BUF1S $T=328600 951000 0 0 $X=328600 $Y=950620
X588 1868 1 2 2052 BUF1S $T=330460 920760 0 0 $X=330460 $Y=920380
X589 117 1 2 138 BUF1S $T=332320 1082040 1 0 $X=332320 $Y=1076620
X590 1920 1 2 2020 BUF1S $T=334180 940920 0 0 $X=334180 $Y=940540
X591 150 1 2 1799 BUF1S $T=343480 1001400 0 180 $X=341000 $Y=995980
X592 1903 1 2 2149 BUF1S $T=344720 1001400 1 0 $X=344720 $Y=995980
X593 129 1 2 157 BUF1S $T=345340 1001400 0 0 $X=345340 $Y=1001020
X594 2149 1 2 2151 BUF1S $T=345340 1051800 1 0 $X=345340 $Y=1046380
X595 99 1 2 160 BUF1S $T=346580 930840 1 0 $X=346580 $Y=925420
X596 162 1 2 1939 BUF1S $T=350920 1011480 0 180 $X=348440 $Y=1006060
X597 168 1 2 2184 BUF1S $T=355880 1082040 1 0 $X=355880 $Y=1076620
X598 119 1 2 164 BUF1S $T=358980 1021560 1 180 $X=356500 $Y=1021180
X599 1790 1 2 174 BUF1S $T=357120 940920 1 0 $X=357120 $Y=935500
X600 2284 1 2 1935 BUF1S $T=367040 1011480 0 180 $X=364560 $Y=1006060
X601 72 1 2 183 BUF1S $T=364560 1082040 0 0 $X=364560 $Y=1081660
X602 195 1 2 182 BUF1S $T=379440 900600 1 180 $X=376960 $Y=900220
X603 2275 1 2 2334 BUF1S $T=378200 1051800 0 0 $X=378200 $Y=1051420
X604 194 1 2 2215 BUF1S $T=380060 900600 0 0 $X=380060 $Y=900220
X605 201 1 2 2248 BUF1S $T=383780 910680 0 180 $X=381300 $Y=905260
X606 202 1 2 1887 BUF1S $T=385020 900600 1 180 $X=382540 $Y=900220
X607 206 1 2 97 BUF1S $T=387500 900600 0 0 $X=387500 $Y=900220
X608 211 1 2 2446 BUF1S $T=391220 1082040 1 0 $X=391220 $Y=1076620
X609 2454 1 2 193 BUF1S $T=403620 1071960 0 180 $X=401140 $Y=1066540
X610 2549 1 2 2398 BUF1S $T=409200 1041720 1 180 $X=406720 $Y=1041340
X611 2601 1 2 2445 BUF1S $T=420980 1021560 0 180 $X=418500 $Y=1016140
X612 2619 1 2 240 BUF1S $T=419120 1051800 1 0 $X=419120 $Y=1046380
X613 2644 1 2 2492 BUF1S $T=424080 1021560 0 180 $X=421600 $Y=1016140
X614 2645 1 2 2465 BUF1S $T=424080 1031640 1 180 $X=421600 $Y=1031260
X615 2650 1 2 2513 BUF1S $T=425320 961080 0 180 $X=422840 $Y=955660
X616 2638 1 2 2600 BUF1S $T=422840 971160 1 0 $X=422840 $Y=965740
X617 2651 1 2 2570 BUF1S $T=427180 971160 1 180 $X=424700 $Y=970780
X618 2652 1 2 2666 BUF1S $T=424700 1021560 1 0 $X=424700 $Y=1016140
X619 2675 1 2 2517 BUF1S $T=429040 1001400 0 180 $X=426560 $Y=995980
X620 2682 1 2 2693 BUF1S $T=429660 920760 0 0 $X=429660 $Y=920380
X621 2702 1 2 2488 BUF1S $T=434620 920760 1 180 $X=432140 $Y=920380
X622 2711 1 2 251 BUF1S $T=434620 1011480 0 180 $X=432140 $Y=1006060
X623 2540 1 2 2710 BUF1S $T=433380 1001400 1 0 $X=433380 $Y=995980
X624 2711 1 2 2607 BUF1S $T=438340 981240 1 180 $X=435860 $Y=980860
X625 2734 1 2 2651 BUF1S $T=441440 971160 0 180 $X=438960 $Y=965740
X626 2734 1 2 2644 BUF1S $T=442060 1001400 0 180 $X=439580 $Y=995980
X627 2747 1 2 2679 BUF1S $T=443300 951000 1 180 $X=440820 $Y=950620
X628 2748 1 2 2619 BUF1S $T=443300 991320 1 180 $X=440820 $Y=990940
X629 270 1 2 267 BUF1S $T=446400 900600 0 0 $X=446400 $Y=900220
X630 2768 1 2 2561 BUF1S $T=450740 971160 1 180 $X=448260 $Y=970780
X631 2793 1 2 2634 BUF1S $T=450740 1031640 1 180 $X=448260 $Y=1031260
X632 268 1 2 2454 BUF1S $T=449500 1021560 0 0 $X=449500 $Y=1021180
X633 2807 1 2 263 BUF1S $T=452600 920760 0 180 $X=450120 $Y=915340
X634 2579 1 2 2767 BUF1S $T=453220 971160 1 180 $X=450740 $Y=970780
X635 2812 1 2 2595 BUF1S $T=453840 961080 1 180 $X=451360 $Y=960700
X636 2813 1 2 2564 BUF1S $T=453840 971160 0 180 $X=451360 $Y=965740
X637 2825 1 2 2734 BUF1S $T=453840 981240 0 180 $X=451360 $Y=975820
X638 2810 1 2 2718 BUF1S $T=453840 1011480 0 180 $X=451360 $Y=1006060
X639 2838 1 2 2450 BUF1S $T=455700 981240 1 180 $X=453220 $Y=980860
X640 2624 1 2 2786 BUF1S $T=453220 991320 0 0 $X=453220 $Y=990940
X641 2718 1 2 2522 BUF1S $T=459420 1031640 1 180 $X=456940 $Y=1031260
X642 2812 1 2 2420 BUF1S $T=463140 1021560 1 180 $X=460660 $Y=1021180
X643 2813 1 2 2385 BUF1S $T=467480 1031640 0 180 $X=465000 $Y=1026220
X644 2888 1 2 2582 BUF1S $T=468100 1031640 1 180 $X=465620 $Y=1031260
X645 2744 1 2 2730 BUF1S $T=469340 951000 0 180 $X=466860 $Y=945580
X646 268 1 2 2902 BUF1S $T=469340 920760 0 0 $X=469340 $Y=920380
X647 2875 1 2 2753 BUF1S $T=469340 930840 0 0 $X=469340 $Y=930460
X648 2906 1 2 2805 BUF1S $T=473680 971160 1 180 $X=471200 $Y=970780
X649 2947 1 2 2711 BUF1S $T=475540 991320 0 180 $X=473060 $Y=985900
X650 305 1 2 2951 BUF1S $T=475540 900600 0 0 $X=475540 $Y=900220
X651 2945 1 2 2813 BUF1S $T=478640 971160 0 180 $X=476160 $Y=965740
X652 2876 1 2 2950 BUF1S $T=476160 1051800 1 0 $X=476160 $Y=1046380
X653 2888 1 2 2642 BUF1S $T=478640 1061880 0 180 $X=476160 $Y=1056460
X654 2948 1 2 2812 BUF1S $T=479260 961080 0 180 $X=476780 $Y=955660
X655 2955 1 2 2828 BUF1S $T=479880 1001400 1 180 $X=477400 $Y=1001020
X656 2942 1 2 2810 BUF1S $T=480500 951000 1 180 $X=478020 $Y=950620
X657 2828 1 2 2887 BUF1S $T=478020 1021560 1 0 $X=478020 $Y=1016140
X658 2949 1 2 2892 BUF1S $T=478640 991320 1 0 $X=478640 $Y=985900
X659 2721 1 2 2979 BUF1S $T=479880 1001400 0 0 $X=479880 $Y=1001020
X660 311 1 2 273 BUF1S $T=486080 930840 0 180 $X=483600 $Y=925420
X661 2540 1 2 2984 BUF1S $T=484840 951000 1 0 $X=484840 $Y=945580
X662 2483 1 2 2884 BUF1S $T=489180 940920 1 0 $X=489180 $Y=935500
X663 3037 1 2 299 BUF1S $T=493520 1051800 1 180 $X=491040 $Y=1051420
X664 3005 1 2 292 BUF1S $T=494760 1061880 0 180 $X=492280 $Y=1056460
X665 3069 1 2 2748 BUF1S $T=500340 981240 1 180 $X=497860 $Y=980860
X666 3106 1 2 322 BUF1S $T=507780 1041720 0 180 $X=505300 $Y=1036300
X667 3114 1 2 3037 BUF1S $T=509020 1011480 0 180 $X=506540 $Y=1006060
X668 3121 1 2 3012 BUF1S $T=510260 1031640 1 180 $X=507780 $Y=1031260
X669 3123 1 2 2601 BUF1S $T=510880 1001400 1 180 $X=508400 $Y=1001020
X670 354 1 2 3071 BUF1S $T=514600 1071960 1 180 $X=512120 $Y=1071580
X671 3141 1 2 3005 BUF1S $T=517080 981240 1 180 $X=514600 $Y=980860
X672 3169 1 2 3114 BUF1S $T=519560 981240 1 180 $X=517080 $Y=980860
X673 3115 1 2 3157 BUF1S $T=518940 1021560 1 0 $X=518940 $Y=1016140
X674 3099 1 2 3180 BUF1S $T=520180 930840 1 0 $X=520180 $Y=925420
X675 340 1 2 286 BUF1S $T=523280 910680 0 180 $X=520800 $Y=905260
X676 3180 1 2 3154 BUF1S $T=520800 930840 0 0 $X=520800 $Y=930460
X677 3203 1 2 3182 BUF1S $T=524520 1001400 1 0 $X=524520 $Y=995980
X678 3059 1 2 3203 BUF1S $T=527000 1001400 1 0 $X=527000 $Y=995980
X679 3123 1 2 3219 BUF1S $T=527000 1011480 1 0 $X=527000 $Y=1006060
X680 3222 1 2 3190 BUF1S $T=530100 951000 0 180 $X=527620 $Y=945580
X681 3115 1 2 3232 BUF1S $T=528860 1031640 1 0 $X=528860 $Y=1026220
X682 365 1 2 3101 BUF1S $T=533200 910680 1 0 $X=533200 $Y=905260
X683 3222 1 2 3121 BUF1S $T=536300 951000 0 180 $X=533820 $Y=945580
X684 3240 1 2 3141 BUF1S $T=537540 971160 1 180 $X=535060 $Y=970780
X685 3209 1 2 3259 BUF1S $T=535060 981240 0 0 $X=535060 $Y=980860
X686 3231 1 2 376 BUF1S $T=537540 1061880 0 180 $X=535060 $Y=1056460
X687 3219 1 2 3277 BUF1S $T=536920 1011480 1 0 $X=536920 $Y=1006060
X688 3280 1 2 3209 BUF1S $T=542500 951000 1 180 $X=540020 $Y=950620
X689 3276 1 2 392 BUF1S $T=540640 1051800 0 0 $X=540640 $Y=1051420
X690 3303 1 2 391 BUF1S $T=544360 1061880 0 180 $X=541880 $Y=1056460
X691 3223 1 2 3307 BUF1S $T=542500 971160 0 0 $X=542500 $Y=970780
X692 3333 1 2 3288 BUF1S $T=548080 951000 1 0 $X=548080 $Y=945580
X693 406 1 2 3358 BUF1S $T=550560 900600 0 0 $X=550560 $Y=900220
X694 407 1 2 3364 BUF1S $T=554900 951000 0 0 $X=554900 $Y=950620
X695 3176 1 2 3399 BUF1S $T=558000 1031640 0 0 $X=558000 $Y=1031260
X696 3321 1 2 3409 BUF1S $T=564200 991320 1 180 $X=561720 $Y=990940
X697 3307 1 2 3407 BUF1S $T=562340 961080 1 0 $X=562340 $Y=955660
X698 3437 1 2 3283 BUF1S $T=567300 1001400 0 180 $X=564820 $Y=995980
X699 3440 1 2 3373 BUF1S $T=567920 971160 0 180 $X=565440 $Y=965740
X700 384 1 2 3437 BUF1S $T=567300 1001400 1 0 $X=567300 $Y=995980
X701 3306 1 2 3391 BUF1S $T=567300 1051800 0 0 $X=567300 $Y=1051420
X702 3440 1 2 3231 BUF1S $T=571020 1011480 0 180 $X=568540 $Y=1006060
X703 3443 1 2 3291 BUF1S $T=571640 1021560 0 180 $X=569160 $Y=1016140
X704 3113 1 2 3464 BUF1S $T=571020 961080 1 0 $X=571020 $Y=955660
X705 3397 1 2 3461 BUF1S $T=574120 920760 1 0 $X=574120 $Y=915340
X706 3271 1 2 3311 BUF1S $T=579700 1001400 0 180 $X=577220 $Y=995980
X707 3496 1 2 3353 BUF1S $T=579700 1021560 0 180 $X=577220 $Y=1016140
X708 3391 1 2 3356 BUF1S $T=577220 1051800 0 0 $X=577220 $Y=1051420
X709 451 1 2 3293 BUF1S $T=577840 951000 1 0 $X=577840 $Y=945580
X710 3306 1 2 3385 BUF1S $T=577840 1031640 1 0 $X=577840 $Y=1026220
X711 3414 1 2 3368 BUF1S $T=582800 951000 0 180 $X=580320 $Y=945580
X712 3385 1 2 3473 BUF1S $T=583420 1011480 1 180 $X=580940 $Y=1011100
X713 3516 1 2 3354 BUF1S $T=584040 1041720 0 180 $X=581560 $Y=1036300
X714 3397 1 2 3511 BUF1S $T=582800 930840 1 0 $X=582800 $Y=925420
X715 3496 1 2 431 BUF1S $T=585280 1041720 1 180 $X=582800 $Y=1041340
X716 3516 1 2 3369 BUF1S $T=583420 1001400 1 0 $X=583420 $Y=995980
X717 3500 1 2 3519 BUF1S $T=589000 961080 0 180 $X=586520 $Y=955660
X718 3385 1 2 3539 BUF1S $T=587140 1011480 1 0 $X=587140 $Y=1006060
X719 3500 1 2 469 BUF1S $T=590240 940920 0 0 $X=590240 $Y=940540
X720 3378 1 2 3417 BUF1S $T=592720 1041720 0 180 $X=590240 $Y=1036300
X721 3558 1 2 3516 BUF1S $T=596440 1001400 0 180 $X=593960 $Y=995980
X722 3586 1 2 3378 BUF1S $T=599540 981240 1 180 $X=597060 $Y=980860
X723 459 1 2 3592 BUF1S $T=598920 1071960 1 0 $X=598920 $Y=1066540
X724 3587 1 2 3023 BUF1S $T=602020 1011480 1 180 $X=599540 $Y=1011100
X725 3582 1 2 3610 BUF1S $T=602020 1011480 0 0 $X=602020 $Y=1011100
X726 3492 1 2 517 BUF1S $T=611940 910680 1 0 $X=611940 $Y=905260
X727 523 1 2 527 BUF1S $T=618140 1082040 0 0 $X=618140 $Y=1081660
X728 3359 1 2 3708 BUF1S $T=618760 951000 1 0 $X=618760 $Y=945580
X729 3657 1 2 502 BUF1S $T=626820 1082040 0 180 $X=624340 $Y=1076620
X730 529 1 2 3676 BUF1S $T=629300 951000 1 180 $X=626820 $Y=950620
X731 3702 1 2 498 BUF1S $T=629920 1082040 1 180 $X=627440 $Y=1081660
X732 3730 1 2 3759 BUF1S $T=631780 1041720 0 180 $X=629300 $Y=1036300
X733 3710 1 2 3794 BUF1S $T=634260 981240 0 0 $X=634260 $Y=980860
X734 3752 1 2 546 BUF1S $T=636120 940920 0 0 $X=636120 $Y=940540
X735 3276 1 2 3806 BUF1S $T=636120 1051800 0 0 $X=636120 $Y=1051420
X736 3812 1 2 3726 BUF1S $T=640460 951000 1 180 $X=637980 $Y=950620
X737 3795 1 2 3657 BUF1S $T=640460 961080 1 180 $X=637980 $Y=960700
X738 3821 1 2 3723 BUF1S $T=642320 930840 1 180 $X=639840 $Y=930460
X739 3834 1 2 3815 BUF1S $T=645420 971160 1 180 $X=642940 $Y=970780
X740 3821 1 2 3669 BUF1S $T=646040 951000 0 180 $X=643560 $Y=945580
X741 3813 1 2 3647 BUF1S $T=646040 1021560 0 180 $X=643560 $Y=1016140
X742 527 1 2 554 BUF1S $T=645420 1082040 0 0 $X=645420 $Y=1081660
X743 3830 1 2 3702 BUF1S $T=648520 971160 1 180 $X=646040 $Y=970780
X744 3858 1 2 3679 BUF1S $T=649760 1001400 0 180 $X=647280 $Y=995980
X745 3860 1 2 3704 BUF1S $T=649760 1011480 0 180 $X=647280 $Y=1006060
X746 3730 1 2 3874 BUF1S $T=650380 1021560 1 0 $X=650380 $Y=1016140
X747 3891 1 2 507 BUF1S $T=655960 1071960 1 180 $X=653480 $Y=1071580
X748 3903 1 2 3821 BUF1S $T=656580 930840 0 180 $X=654100 $Y=925420
X749 3883 1 2 3895 BUF1S $T=654100 940920 0 0 $X=654100 $Y=940540
X750 3891 1 2 3754 BUF1S $T=655340 971160 1 0 $X=655340 $Y=965740
X751 3860 1 2 3644 BUF1S $T=657820 1051800 0 180 $X=655340 $Y=1046380
X752 3858 1 2 3684 BUF1S $T=655960 1031640 0 0 $X=655960 $Y=1031260
X753 3903 1 2 593 BUF1S $T=657820 920760 1 0 $X=657820 $Y=915340
X754 587 1 2 3778 BUF1S $T=659680 951000 1 0 $X=659680 $Y=945580
X755 3940 1 2 3830 BUF1S $T=663400 981240 0 180 $X=660920 $Y=975820
X756 3938 1 2 3682 BUF1S $T=664020 1041720 1 180 $X=661540 $Y=1041340
X757 3813 1 2 3938 BUF1S $T=662160 1011480 0 0 $X=662160 $Y=1011100
X758 3812 1 2 597 BUF1S $T=664020 1082040 0 0 $X=664020 $Y=1081660
X759 601 1 2 3741 BUF1S $T=668980 971160 0 180 $X=666500 $Y=965740
X760 3994 1 2 3085 BUF1S $T=671460 961080 0 180 $X=668980 $Y=955660
X761 3975 1 2 605 BUF1S $T=670220 940920 0 0 $X=670220 $Y=940540
X762 4008 1 2 3748 BUF1S $T=674560 981240 1 180 $X=672080 $Y=980860
X763 3972 1 2 3890 BUF1S $T=672080 1071960 1 0 $X=672080 $Y=1066540
X764 3890 1 2 4019 BUF1S $T=673940 1061880 0 0 $X=673940 $Y=1061500
X765 4019 1 2 612 BUF1S $T=676420 1082040 0 180 $X=673940 $Y=1076620
X766 4029 1 2 3758 BUF1S $T=677660 991320 0 180 $X=675180 $Y=985900
X767 4024 1 2 3901 BUF1S $T=677660 991320 1 180 $X=675180 $Y=990940
X768 3922 1 2 3917 BUF1S $T=676420 981240 1 0 $X=676420 $Y=975820
X769 557 1 2 3587 BUF1S $T=680140 1011480 0 0 $X=680140 $Y=1011100
X770 587 1 2 633 BUF1S $T=682000 1082040 0 0 $X=682000 $Y=1081660
X771 4078 1 2 3774 BUF1S $T=685100 1011480 0 180 $X=682620 $Y=1006060
X772 4100 1 2 3757 BUF1S $T=689440 1011480 1 180 $X=686960 $Y=1011100
X773 605 1 2 644 BUF1S $T=688200 1082040 0 0 $X=688200 $Y=1081660
X774 4000 1 2 4036 BUF1S $T=688820 1001400 1 0 $X=688820 $Y=995980
X775 4108 1 2 4123 BUF1S $T=690680 981240 1 0 $X=690680 $Y=975820
X776 4153 1 2 4003 BUF1S $T=695640 940920 0 180 $X=693160 $Y=935500
X777 4120 1 2 4117 BUF1S $T=694400 1061880 0 0 $X=694400 $Y=1061500
X778 4164 1 2 4088 BUF1S $T=700600 961080 0 180 $X=698120 $Y=955660
X779 4064 1 2 4058 BUF1S $T=700600 971160 0 180 $X=698120 $Y=965740
X780 4087 1 2 4151 BUF1S $T=700600 961080 0 0 $X=700600 $Y=960700
X781 4088 1 2 655 BUF1S $T=700600 1071960 0 0 $X=700600 $Y=1071580
X782 4171 1 2 4086 BUF1S $T=706180 1011480 0 180 $X=703700 $Y=1006060
X783 4164 1 2 4192 BUF1S $T=704940 951000 0 0 $X=704940 $Y=950620
X784 4151 1 2 648 BUF1S $T=705560 1071960 0 0 $X=705560 $Y=1071580
X785 4211 1 2 4216 BUF1S $T=706800 961080 1 0 $X=706800 $Y=955660
X786 4227 1 2 4080 BUF1S $T=709900 940920 1 180 $X=707420 $Y=940540
X787 3846 1 2 4193 BUF1S $T=707420 991320 1 0 $X=707420 $Y=985900
X788 4197 1 2 4176 BUF1S $T=709280 971160 0 0 $X=709280 $Y=970780
X789 630 1 2 4247 BUF1S $T=711140 1071960 0 0 $X=711140 $Y=1071580
X790 4236 1 2 4124 BUF1S $T=713000 1051800 1 0 $X=713000 $Y=1046380
X791 4217 1 2 4253 BUF1S $T=714240 1001400 1 0 $X=714240 $Y=995980
X792 4238 1 2 4259 BUF1S $T=719200 1011480 1 0 $X=719200 $Y=1006060
X793 4253 1 2 4248 BUF1S $T=719820 981240 1 0 $X=719820 $Y=975820
X794 4291 1 2 4066 BUF1S $T=724160 1001400 0 180 $X=721680 $Y=995980
X795 4308 1 2 4061 BUF1S $T=726640 1051800 0 0 $X=726640 $Y=1051420
X796 4221 1 2 4268 BUF1S $T=727260 1061880 0 0 $X=727260 $Y=1061500
X797 676 1 2 4005 BUF1S $T=730360 951000 1 0 $X=730360 $Y=945580
X798 4365 1 2 4001 BUF1S $T=734080 951000 1 180 $X=731600 $Y=950620
X799 4287 1 2 4312 BUF1S $T=732840 920760 0 0 $X=732840 $Y=920380
X800 4227 1 2 701 BUF1S $T=738420 940920 1 180 $X=735940 $Y=940540
X801 4335 1 2 4402 BUF1S $T=738420 920760 1 0 $X=738420 $Y=915340
X802 4332 1 2 4405 BUF1S $T=741520 961080 1 0 $X=741520 $Y=955660
X803 4282 1 2 4403 BUF1S $T=744000 961080 1 0 $X=744000 $Y=955660
X804 717 1 2 675 BUF1S $T=747100 900600 1 180 $X=744620 $Y=900220
X805 718 1 2 4015 BUF1S $T=748960 961080 0 180 $X=746480 $Y=955660
X806 720 1 2 4263 BUF1S $T=750200 930840 0 0 $X=750200 $Y=930460
X807 4463 1 2 4434 BUF1S $T=752680 930840 0 0 $X=752680 $Y=930460
X808 4482 1 2 4401 BUF1S $T=757640 1041720 1 180 $X=755160 $Y=1041340
X809 4486 1 2 4497 BUF1S $T=758260 951000 1 0 $X=758260 $Y=945580
X810 4504 1 2 4452 BUF1S $T=760740 940920 1 0 $X=760740 $Y=935500
X811 4461 1 2 4518 BUF1S $T=760740 940920 0 0 $X=760740 $Y=940540
X812 4522 1 2 727 BUF1S $T=764460 1071960 0 180 $X=761980 $Y=1066540
X813 4523 1 2 4513 BUF1S $T=766940 1041720 0 180 $X=764460 $Y=1036300
X814 4513 1 2 732 BUF1S $T=764460 1071960 1 0 $X=764460 $Y=1066540
X815 4466 1 2 4476 BUF1S $T=765700 951000 0 0 $X=765700 $Y=950620
X816 4539 1 2 4505 BUF1S $T=768180 971160 1 180 $X=765700 $Y=970780
X817 4525 1 2 4455 BUF1S $T=766320 971160 1 0 $X=766320 $Y=965740
X818 4526 1 2 4382 BUF1S $T=769420 1011480 0 0 $X=769420 $Y=1011100
X819 4498 1 2 4553 BUF1S $T=770040 910680 1 0 $X=770040 $Y=905260
X820 4569 1 2 4603 BUF1S $T=771280 920760 0 0 $X=771280 $Y=920380
X821 4539 1 2 4547 BUF1S $T=771280 940920 0 0 $X=771280 $Y=940540
X822 4579 1 2 4557 BUF1S $T=773760 1031640 1 180 $X=771280 $Y=1031260
X823 4146 1 2 4578 BUF1S $T=773140 940920 1 0 $X=773140 $Y=935500
X824 754 1 2 4565 BUF1S $T=775620 1061880 1 180 $X=773140 $Y=1061500
X825 4516 1 2 4485 BUF1S $T=773760 1031640 0 0 $X=773760 $Y=1031260
X826 731 1 2 4604 BUF1S $T=773760 1071960 0 0 $X=773760 $Y=1071580
X827 4593 1 2 4523 BUF1S $T=777480 1021560 0 180 $X=775000 $Y=1016140
X828 4606 1 2 4544 BUF1S $T=776860 1031640 0 0 $X=776860 $Y=1031260
X829 4365 1 2 4568 BUF1S $T=777480 1021560 1 0 $X=777480 $Y=1016140
X830 4618 1 2 4599 BUF1S $T=778720 1011480 1 0 $X=778720 $Y=1006060
X831 4580 1 2 4636 BUF1S $T=779340 1051800 0 0 $X=779340 $Y=1051420
X832 4654 1 2 4577 BUF1S $T=784920 930840 1 0 $X=784920 $Y=925420
X833 4656 1 2 4668 BUF1S $T=784920 1021560 0 0 $X=784920 $Y=1021180
X834 4005 1 2 4639 BUF1S $T=787400 1021560 0 0 $X=787400 $Y=1021180
X835 4692 1 2 4620 BUF1S $T=791740 940920 1 180 $X=789260 $Y=940540
X836 4695 1 2 4637 BUF1S $T=791740 971160 0 180 $X=789260 $Y=965740
X837 4692 1 2 4719 BUF1S $T=790500 940920 1 0 $X=790500 $Y=935500
X838 4482 1 2 4708 BUF1S $T=791120 1051800 0 0 $X=791120 $Y=1051420
X839 4709 1 2 788 BUF1S $T=793600 1071960 1 180 $X=791120 $Y=1071580
X840 4734 1 2 4742 BUF1S $T=795460 1011480 0 0 $X=795460 $Y=1011100
X841 808 1 2 4757 BUF1S $T=797320 900600 0 0 $X=797320 $Y=900220
X842 620 1 2 4761 BUF1S $T=799800 930840 1 0 $X=799800 $Y=925420
X843 4775 1 2 4709 BUF1S $T=802280 1041720 1 180 $X=799800 $Y=1041340
X844 4803 1 2 4729 BUF1S $T=806620 961080 1 180 $X=804140 $Y=960700
X845 4813 1 2 4718 BUF1S $T=807860 971160 1 180 $X=805380 $Y=970780
X846 4861 1 2 779 BUF1S $T=816540 910680 1 180 $X=814060 $Y=910300
X847 4853 1 2 4884 BUF1S $T=816540 1041720 0 0 $X=816540 $Y=1041340
X848 4884 1 2 821 BUF1S $T=819020 1071960 1 0 $X=819020 $Y=1066540
X849 4903 1 2 4910 BUF1S $T=820880 1011480 0 0 $X=820880 $Y=1011100
X850 4859 1 2 4881 BUF1S $T=822120 1061880 1 0 $X=822120 $Y=1056460
X851 4904 1 2 4763 BUF1S $T=822740 1021560 0 0 $X=822740 $Y=1021180
X852 346 1 2 4896 BUF1S $T=823980 961080 1 0 $X=823980 $Y=955660
X853 841 1 2 850 BUF1S $T=823980 1082040 1 0 $X=823980 $Y=1076620
X854 805 1 2 851 BUF1S $T=827080 910680 1 180 $X=824600 $Y=910300
X855 803 1 2 4933 BUF1S $T=826460 910680 1 0 $X=826460 $Y=905260
X856 4923 1 2 818 BUF1S $T=828940 1082040 0 180 $X=826460 $Y=1076620
X857 4886 1 2 4944 BUF1S $T=827080 1001400 0 0 $X=827080 $Y=1001020
X858 4908 1 2 4914 BUF1S $T=828940 940920 1 0 $X=828940 $Y=935500
X859 4872 1 2 4923 BUF1S $T=828940 1041720 0 0 $X=828940 $Y=1041340
X860 789 1 2 4959 BUF1S $T=831420 910680 1 0 $X=831420 $Y=905260
X861 4114 1 2 4955 BUF1S $T=832040 920760 0 0 $X=832040 $Y=920380
X862 4977 1 2 864 BUF1S $T=837620 1082040 0 180 $X=835140 $Y=1076620
X863 4951 1 2 4856 BUF1S $T=840100 1041720 1 180 $X=837620 $Y=1041340
X864 4883 1 2 4995 BUF1S $T=838860 910680 0 0 $X=838860 $Y=910300
X865 842 1 2 4966 BUF1S $T=838860 940920 1 0 $X=838860 $Y=935500
X866 5007 1 2 4977 BUF1S $T=842580 1021560 1 180 $X=840100 $Y=1021180
X867 350 1 2 5020 BUF1S $T=841960 930840 0 0 $X=841960 $Y=930460
X868 4609 1 2 5018 BUF1S $T=844440 940920 0 0 $X=844440 $Y=940540
X869 861 1 2 862 BUF1S $T=844440 1082040 0 0 $X=844440 $Y=1081660
X870 4797 1 2 5054 BUF1S $T=847540 1041720 1 0 $X=847540 $Y=1036300
X871 5031 1 2 5063 BUF1S $T=851260 1031640 1 0 $X=851260 $Y=1026220
X872 5072 1 2 5079 BUF1S $T=852500 1031640 0 0 $X=852500 $Y=1031260
X873 5055 1 2 5101 BUF1S $T=853120 1011480 0 0 $X=853120 $Y=1011100
X874 5078 1 2 5085 BUF1S $T=856840 920760 1 0 $X=856840 $Y=915340
X875 5108 1 2 4961 BUF1S $T=859320 951000 0 180 $X=856840 $Y=945580
X876 4961 1 2 5109 BUF1S $T=856840 961080 0 0 $X=856840 $Y=960700
X877 4952 1 2 5114 BUF1S $T=858080 991320 0 0 $X=858080 $Y=990940
X878 5095 1 2 880 BUF1S $T=861180 1071960 0 180 $X=858700 $Y=1066540
X879 4992 1 2 5124 BUF1S $T=859320 961080 0 0 $X=859320 $Y=960700
X880 5032 1 2 5095 BUF1S $T=861180 1021560 0 0 $X=861180 $Y=1021180
X881 4997 1 2 5147 BUF1S $T=861800 961080 0 0 $X=861800 $Y=960700
X882 862 1 2 5143 BUF1S $T=863040 1051800 1 0 $X=863040 $Y=1046380
X883 5140 1 2 5067 BUF1S $T=868000 951000 1 180 $X=865520 $Y=950620
X884 5083 1 2 5179 BUF1S $T=868620 920760 1 0 $X=868620 $Y=915340
X885 4967 1 2 5138 BUF1S $T=868620 951000 1 0 $X=868620 $Y=945580
X886 5149 1 2 909 BUF1S $T=873580 1071960 1 0 $X=873580 $Y=1066540
X887 4997 1 2 5225 BUF1S $T=876060 951000 0 0 $X=876060 $Y=950620
X888 4992 1 2 5242 BUF1S $T=878540 951000 0 0 $X=878540 $Y=950620
X889 5196 1 2 5140 BUF1S $T=881020 961080 1 180 $X=878540 $Y=960700
X890 4967 1 2 5255 BUF1S $T=879780 940920 0 0 $X=879780 $Y=940540
X891 923 1 2 5248 BUF1S $T=882880 1071960 0 180 $X=880400 $Y=1066540
X892 5108 1 2 5277 BUF1S $T=882880 940920 0 0 $X=882880 $Y=940540
X893 5114 1 2 5284 BUF1S $T=884740 991320 1 0 $X=884740 $Y=985900
X894 5196 1 2 5287 BUF1S $T=885360 971160 0 0 $X=885360 $Y=970780
X895 5143 1 2 5265 BUF1S $T=887840 1051800 0 180 $X=885360 $Y=1046380
X896 5298 1 2 5306 BUF1S $T=887220 1061880 1 0 $X=887220 $Y=1056460
X897 5021 1 2 5338 BUF1S $T=890320 991320 1 0 $X=890320 $Y=985900
X898 5213 1 2 5300 BUF1S $T=890320 1041720 1 0 $X=890320 $Y=1036300
X899 5213 1 2 917 BUF1S $T=892800 1071960 0 180 $X=890320 $Y=1066540
X900 5245 1 2 941 BUF1S $T=892800 1071960 1 0 $X=892800 $Y=1066540
X901 5287 1 2 5340 BUF1S $T=896520 981240 0 0 $X=896520 $Y=980860
X902 5268 1 2 5352 BUF1S $T=897760 1001400 0 0 $X=897760 $Y=1001020
X903 5284 1 2 5372 BUF1S $T=899000 991320 0 0 $X=899000 $Y=990940
X904 5204 1 2 5333 BUF1S $T=902720 1021560 0 0 $X=902720 $Y=1021180
X905 5320 1 2 5313 BUF1S $T=903960 1031640 0 0 $X=903960 $Y=1031260
X906 5399 1 2 5321 BUF1S $T=908920 930840 0 180 $X=906440 $Y=925420
X907 938 1 2 5406 BUF1S $T=908300 1071960 0 0 $X=908300 $Y=1071580
X908 5263 1 2 5415 BUF1S $T=913880 981240 0 0 $X=913880 $Y=980860
X909 5399 1 2 5446 BUF1S $T=918220 920760 0 0 $X=918220 $Y=920380
X910 958 1 2 5223 BUF1S $T=920700 951000 0 180 $X=918220 $Y=945580
X911 5458 1 2 5476 BUF1S $T=921320 961080 0 0 $X=921320 $Y=960700
X912 993 1 2 5463 BUF1S $T=926280 940920 0 180 $X=923800 $Y=935500
X913 5523 1 2 5442 BUF1S $T=931860 1031640 1 180 $X=929380 $Y=1031260
X914 987 1 2 5498 BUF1S $T=930000 920760 0 0 $X=930000 $Y=920380
X915 5490 1 2 5527 BUF1S $T=930000 961080 0 0 $X=930000 $Y=960700
X916 5537 1 2 5523 BUF1S $T=935580 971160 1 180 $X=933100 $Y=970780
X917 5527 1 2 991 BUF1S $T=933100 1082040 0 0 $X=933100 $Y=1081660
X918 3962 1 2 5577 BUF1S $T=937440 961080 0 0 $X=937440 $Y=960700
X919 5559 1 2 5453 BUF1S $T=939920 1041720 1 180 $X=937440 $Y=1041340
X920 5487 1 2 5589 BUF1S $T=938060 971160 0 0 $X=938060 $Y=970780
X921 5562 1 2 972 BUF1S $T=938680 1082040 0 0 $X=938680 $Y=1081660
X922 5457 1 2 5562 BUF1S $T=941780 971160 0 0 $X=941780 $Y=970780
X923 5592 1 2 5550 BUF1S $T=942400 981240 1 0 $X=942400 $Y=975820
X924 5526 1 2 5636 BUF1S $T=947360 951000 0 0 $X=947360 $Y=950620
X925 5529 1 2 5650 BUF1S $T=947980 1021560 1 0 $X=947980 $Y=1016140
X926 5626 1 2 5643 BUF1S $T=947980 1031640 1 0 $X=947980 $Y=1026220
X927 5262 1 2 1026 BUF1S $T=951700 1082040 0 180 $X=949220 $Y=1076620
X928 5576 1 2 5618 BUF1S $T=952320 920760 0 0 $X=952320 $Y=920380
X929 1028 1 2 5654 BUF1S $T=952320 991320 1 0 $X=952320 $Y=985900
X930 1031 1 2 5646 BUF1S $T=952940 1011480 0 0 $X=952940 $Y=1011100
X931 1007 1 2 1035 BUF1S $T=954180 900600 0 0 $X=954180 $Y=900220
X932 5610 1 2 5678 BUF1S $T=959140 971160 1 180 $X=956660 $Y=970780
X933 5631 1 2 5704 BUF1S $T=957280 910680 0 0 $X=957280 $Y=910300
X934 5685 1 2 5696 BUF1S $T=957900 991320 0 0 $X=957900 $Y=990940
X935 5678 1 2 1036 BUF1S $T=960380 1071960 0 180 $X=957900 $Y=1066540
X936 1028 1 2 5687 BUF1S $T=959140 951000 0 0 $X=959140 $Y=950620
X937 1021 1 2 5707 BUF1S $T=959760 940920 1 0 $X=959760 $Y=935500
X938 5721 1 2 1050 BUF1S $T=965340 1071960 0 180 $X=962860 $Y=1066540
X939 5717 1 2 5532 BUF1S $T=967200 1021560 1 180 $X=964720 $Y=1021180
X940 5682 1 2 5652 BUF1S $T=966580 920760 0 0 $X=966580 $Y=920380
X941 5603 1 2 5721 BUF1S $T=971540 971160 0 180 $X=969060 $Y=965740
X942 5743 1 2 5560 BUF1S $T=971540 1051800 0 180 $X=969060 $Y=1046380
X943 5765 1 2 1023 BUF1S $T=974640 910680 1 180 $X=972160 $Y=910300
X944 5669 1 2 5779 BUF1S $T=972160 961080 0 0 $X=972160 $Y=960700
X945 1052 1 2 5548 BUF1S $T=974020 940920 1 0 $X=974020 $Y=935500
X946 5779 1 2 5657 BUF1S $T=976500 1021560 1 180 $X=974020 $Y=1021180
X947 5796 1 2 5627 BUF1S $T=978360 1031640 1 180 $X=975880 $Y=1031260
X948 5717 1 2 5743 BUF1S $T=977120 1021560 0 0 $X=977120 $Y=1021180
X949 5635 1 2 5796 BUF1S $T=978980 940920 0 0 $X=978980 $Y=940540
X950 5717 1 2 5804 BUF1S $T=979600 1021560 0 0 $X=979600 $Y=1021180
X951 5804 1 2 5719 BUF1S $T=980840 1011480 0 0 $X=980840 $Y=1011100
X952 5763 1 2 1065 BUF1S $T=983940 1071960 1 180 $X=981460 $Y=1071580
X953 5763 1 2 1076 BUF1S $T=984560 1071960 0 0 $X=984560 $Y=1071580
X954 5697 1 2 5732 BUF1S $T=989520 971160 1 180 $X=987040 $Y=970780
X955 5828 1 2 5810 BUF1S $T=988280 940920 0 0 $X=988280 $Y=940540
X956 5810 1 2 5829 BUF1S $T=988280 981240 0 0 $X=988280 $Y=980860
X957 5497 1 2 5757 BUF1S $T=990760 991320 1 180 $X=988280 $Y=990940
X958 5719 1 2 5697 BUF1S $T=990760 1001400 0 180 $X=988280 $Y=995980
X959 5847 1 2 5763 BUF1S $T=992620 1051800 1 180 $X=990140 $Y=1051420
X960 5765 1 2 1078 BUF1S $T=993860 920760 1 180 $X=991380 $Y=920380
X961 5719 1 2 5854 BUF1S $T=991380 991320 0 0 $X=991380 $Y=990940
X962 5829 1 2 1084 BUF1S $T=991380 1031640 0 0 $X=991380 $Y=1031260
X963 5765 1 2 1086 BUF1S $T=993860 910680 0 0 $X=993860 $Y=910300
X964 5865 1 2 5851 BUF1S $T=996340 940920 0 0 $X=996340 $Y=940540
X965 5857 1 2 5867 BUF1S $T=996960 1031640 1 0 $X=996960 $Y=1026220
X966 5887 1 2 5870 BUF1S $T=1001300 1001400 1 180 $X=998820 $Y=1001020
X967 5729 1 2 5900 BUF1S $T=1000060 1031640 1 0 $X=1000060 $Y=1026220
X968 5883 1 2 5903 BUF1S $T=1000680 981240 1 0 $X=1000680 $Y=975820
X969 5905 1 2 5915 BUF1S $T=1003780 940920 0 0 $X=1003780 $Y=940540
X970 5847 1 2 5910 BUF1S $T=1003780 1051800 1 0 $X=1003780 $Y=1046380
X971 5897 1 2 1108 BUF1S $T=1004400 1041720 1 0 $X=1004400 $Y=1036300
X972 5854 1 2 5872 BUF1S $T=1009360 981240 1 0 $X=1009360 $Y=975820
X973 5962 1 2 5920 BUF1S $T=1013080 940920 1 0 $X=1013080 $Y=935500
X974 1116 1 2 5962 BUF1S $T=1013080 940920 0 0 $X=1013080 $Y=940540
X975 5915 1 2 5986 BUF1S $T=1014940 981240 1 0 $X=1014940 $Y=975820
X976 5986 1 2 1129 BUF1S $T=1017420 1041720 0 180 $X=1014940 $Y=1036300
X977 5968 1 2 5901 BUF1S $T=1016180 910680 0 0 $X=1016180 $Y=910300
X978 958 1 2 5852 BUF1S $T=1016180 940920 0 0 $X=1016180 $Y=940540
X979 1132 1 2 5961 BUF1S $T=1016800 920760 1 0 $X=1016800 $Y=915340
X980 6000 1 2 6026 BUF1S $T=1021760 951000 1 0 $X=1021760 $Y=945580
X981 6026 1 2 6027 BUF1S $T=1023620 991320 1 0 $X=1023620 $Y=985900
X982 5938 1 2 6018 BUF1S $T=1025480 920760 0 0 $X=1025480 $Y=920380
X983 6027 1 2 1151 BUF1S $T=1031060 1041720 1 180 $X=1028580 $Y=1041340
X984 6073 1 2 6083 BUF1S $T=1031680 1051800 1 0 $X=1031680 $Y=1046380
X985 5852 1 2 6071 BUF1S $T=1033540 940920 0 0 $X=1033540 $Y=940540
X986 6081 1 2 6091 BUF1S $T=1033540 971160 1 0 $X=1033540 $Y=965740
X987 6079 1 2 6092 BUF1S $T=1033540 1041720 1 0 $X=1033540 $Y=1036300
X988 1158 1 2 6096 BUF1S $T=1034160 910680 0 0 $X=1034160 $Y=910300
X989 5994 1 2 6070 BUF1S $T=1034780 910680 1 0 $X=1034780 $Y=905260
X990 6080 1 2 1156 BUF1S $T=1036020 1041720 1 0 $X=1036020 $Y=1036300
X991 6116 1 2 1160 BUF1S $T=1040360 1031640 1 180 $X=1037880 $Y=1031260
X992 6091 1 2 6116 BUF1S $T=1039740 991320 0 0 $X=1039740 $Y=990940
X993 1166 1 2 6028 BUF1S $T=1040360 910680 1 0 $X=1040360 $Y=905260
X994 6119 1 2 6142 BUF1S $T=1042840 971160 1 0 $X=1042840 $Y=965740
X995 5968 1 2 6153 BUF1S $T=1044700 910680 0 0 $X=1044700 $Y=910300
X996 6125 1 2 6145 BUF1S $T=1045940 940920 1 0 $X=1045940 $Y=935500
X997 6162 1 2 6029 BUF1S $T=1049040 951000 1 180 $X=1046560 $Y=950620
X998 6088 1 2 6168 BUF1S $T=1048420 940920 1 0 $X=1048420 $Y=935500
X999 1161 1 2 1187 BUF1S $T=1049660 900600 0 0 $X=1049660 $Y=900220
X1000 6192 1 2 6191 BUF1S $T=1055860 940920 0 0 $X=1055860 $Y=940540
X1001 6064 1 2 6099 BUF1S $T=1056480 971160 0 0 $X=1056480 $Y=970780
X1002 6093 1 2 6187 BUF1S $T=1057100 1031640 0 0 $X=1057100 $Y=1031260
X1003 6144 1 2 6194 BUF1S $T=1058960 1021560 0 0 $X=1058960 $Y=1021180
X1004 6232 1 2 6148 BUF1S $T=1062680 951000 0 0 $X=1062680 $Y=950620
X1005 1161 1 2 6167 BUF1S $T=1067020 920760 1 180 $X=1064540 $Y=920380
X1006 6259 1 2 6126 BUF1S $T=1068260 1001400 0 180 $X=1065780 $Y=995980
X1007 6277 1 2 6169 BUF1S $T=1071360 1001400 0 0 $X=1071360 $Y=1001020
X1008 6290 1 2 6240 BUF1S $T=1075700 1011480 0 180 $X=1073220 $Y=1006060
X1009 6159 1 2 6295 BUF1S $T=1075080 910680 1 0 $X=1075080 $Y=905260
X1010 6231 1 2 6202 BUF1S $T=1077560 971160 0 180 $X=1075080 $Y=965740
X1011 6146 1 2 6312 BUF1S $T=1076940 940920 1 0 $X=1076940 $Y=935500
X1012 6303 1 2 6265 BUF1S $T=1079420 1011480 0 180 $X=1076940 $Y=1006060
X1013 6236 1 2 6333 BUF1S $T=1081900 1051800 1 0 $X=1081900 $Y=1046380
X1014 6277 1 2 6338 BUF1S $T=1081900 1071960 1 0 $X=1081900 $Y=1066540
X1015 6168 1 2 6290 BUF1S $T=1085000 951000 1 180 $X=1082520 $Y=950620
X1016 6192 1 2 6321 BUF1S $T=1082520 1061880 0 0 $X=1082520 $Y=1061500
X1017 6145 1 2 6303 BUF1S $T=1083760 951000 1 0 $X=1083760 $Y=945580
X1018 6259 1 2 6346 BUF1S $T=1084380 1001400 0 0 $X=1084380 $Y=1001020
X1019 6359 1 2 1234 BUF1S $T=1089960 1001400 1 180 $X=1087480 $Y=1001020
X1020 6197 1 2 6370 BUF1S $T=1093680 930840 1 0 $X=1093680 $Y=925420
X1021 1247 1 2 6199 BUF1S $T=1096160 961080 1 180 $X=1093680 $Y=960700
X1022 6370 1 2 1230 BUF1S $T=1093680 1011480 1 0 $X=1093680 $Y=1006060
X1023 6186 1 2 6359 BUF1S $T=1096160 930840 1 0 $X=1096160 $Y=925420
X1024 6190 1 2 6408 BUF1S $T=1096160 961080 0 0 $X=1096160 $Y=960700
X1025 6167 1 2 6332 BUF1S $T=1098640 930840 1 0 $X=1098640 $Y=925420
X1026 6181 1 2 6415 BUF1S $T=1098640 951000 1 0 $X=1098640 $Y=945580
X1027 6363 1 2 6398 BUF1S $T=1099880 961080 0 0 $X=1099880 $Y=960700
X1028 6287 1 2 6440 BUF1S $T=1103600 961080 0 0 $X=1103600 $Y=960700
X1029 6408 1 2 1245 BUF1S $T=1106080 1001400 1 180 $X=1103600 $Y=1001020
X1030 6312 1 2 6477 BUF1S $T=1105460 940920 0 0 $X=1105460 $Y=940540
X1031 6447 1 2 6400 BUF1S $T=1106080 1001400 0 0 $X=1106080 $Y=1001020
X1032 6333 1 2 6450 BUF1S $T=1111660 1051800 0 180 $X=1109180 $Y=1046380
X1033 6415 1 2 1268 BUF1S $T=1110420 1011480 1 0 $X=1110420 $Y=1006060
X1034 6421 1 2 6472 BUF1S $T=1112900 1011480 1 0 $X=1112900 $Y=1006060
X1035 6231 1 2 6510 BUF1S $T=1115380 971160 1 0 $X=1115380 $Y=965740
X1036 6333 1 2 6512 BUF1S $T=1115380 1051800 0 0 $X=1115380 $Y=1051420
X1037 6512 1 2 1250 BUF1S $T=1118480 1061880 1 180 $X=1116000 $Y=1061500
X1038 6500 1 2 6492 BUF1S $T=1116620 981240 1 0 $X=1116620 $Y=975820
X1039 1214 1 2 1282 BUF1S $T=1117860 910680 0 0 $X=1117860 $Y=910300
X1040 6255 1 2 6486 BUF1S $T=1117860 991320 0 0 $X=1117860 $Y=990940
X1041 6510 1 2 6441 BUF1S $T=1127780 1011480 1 180 $X=1125300 $Y=1011100
X1042 1338 1 2 1374 DELB $T=226300 981240 1 0 $X=226300 $Y=975820
X1043 1402 1 2 1413 DELB $T=236840 991320 0 0 $X=236840 $Y=990940
X1044 1447 1 2 1463 DELB $T=244280 991320 0 0 $X=244280 $Y=990940
X1045 1554 1 2 1723 DELB $T=277760 991320 0 0 $X=277760 $Y=990940
X1046 1870 1 2 85 DELB $T=303180 1071960 0 0 $X=303180 $Y=1071580
X1047 1952 1 2 114 DELB $T=315580 1082040 1 0 $X=315580 $Y=1076620
X1048 2007 1 2 2034 DELB $T=326120 981240 0 0 $X=326120 $Y=980860
X1049 2129 1 2 2155 DELB $T=342860 1041720 0 0 $X=342860 $Y=1041340
X1050 2109 1 2 2111 DELB $T=345960 1071960 1 0 $X=345960 $Y=1066540
X1051 2175 1 2 2098 DELB $T=350300 1082040 1 0 $X=350300 $Y=1076620
X1052 2182 1 2 2183 DELB $T=351540 1011480 1 0 $X=351540 $Y=1006060
X1053 2194 1 2 2203 DELB $T=352780 1041720 1 0 $X=352780 $Y=1036300
X1054 2222 1 2 2242 DELB $T=357120 981240 1 0 $X=357120 $Y=975820
X1055 2236 1 2 2257 DELB $T=359600 1011480 1 0 $X=359600 $Y=1006060
X1056 2329 1 2 2359 DELB $T=373860 1061880 0 0 $X=373860 $Y=1061500
X1057 2332 1 2 2328 DELB $T=374480 1001400 0 0 $X=374480 $Y=1001020
X1058 2438 1 2 2467 DELB $T=391220 961080 0 0 $X=391220 $Y=960700
X1059 2440 1 2 2470 DELB $T=394940 1082040 1 0 $X=394940 $Y=1076620
X1060 2461 1 2 2474 DELB $T=396800 1021560 0 0 $X=396800 $Y=1021180
X1061 2496 1 2 2524 DELB $T=401140 930840 1 0 $X=401140 $Y=925420
X1062 2526 1 2 2527 DELB $T=405480 1031640 1 0 $X=405480 $Y=1026220
X1063 2528 1 2 2521 DELB $T=405480 1051800 0 0 $X=405480 $Y=1051420
X1064 2548 1 2 2575 DELB $T=408580 951000 0 0 $X=408580 $Y=950620
X1065 2520 1 2 2510 DELB $T=411060 1011480 0 0 $X=411060 $Y=1011100
X1066 2534 1 2 2586 DELB $T=414780 1031640 1 0 $X=414780 $Y=1026220
X1067 2541 1 2 2587 DELB $T=414780 1051800 0 0 $X=414780 $Y=1051420
X1068 2589 1 2 2615 DELB $T=414780 1082040 0 0 $X=414780 $Y=1081660
X1069 2598 1 2 2626 DELB $T=416020 930840 0 0 $X=416020 $Y=930460
X1070 2611 1 2 2657 DELB $T=422220 1031640 1 0 $X=422220 $Y=1026220
X1071 2647 1 2 2670 DELB $T=424080 1071960 1 0 $X=424080 $Y=1066540
X1072 2689 1 2 2713 DELB $T=430900 981240 0 0 $X=430900 $Y=980860
X1073 2722 1 2 2727 DELB $T=435860 951000 0 0 $X=435860 $Y=950620
X1074 2694 1 2 2677 DELB $T=436480 1031640 0 0 $X=436480 $Y=1031260
X1075 2740 1 2 2762 DELB $T=440200 1061880 1 0 $X=440200 $Y=1056460
X1076 2743 1 2 2754 DELB $T=441440 981240 0 0 $X=441440 $Y=980860
X1077 2774 1 2 2780 DELB $T=446400 971160 1 0 $X=446400 $Y=965740
X1078 2705 1 2 2745 DELB $T=446400 1031640 1 0 $X=446400 $Y=1026220
X1079 2776 1 2 2781 DELB $T=448260 981240 0 0 $X=448260 $Y=980860
X1080 2772 1 2 2752 DELB $T=449500 1061880 0 0 $X=449500 $Y=1061500
X1081 2798 1 2 2822 DELB $T=450120 1061880 1 0 $X=450120 $Y=1056460
X1082 2809 1 2 2829 DELB $T=452600 1021560 0 0 $X=452600 $Y=1021180
X1083 2843 1 2 2842 DELB $T=458180 1061880 0 0 $X=458180 $Y=1061500
X1084 2834 1 2 2832 DELB $T=461280 1041720 1 0 $X=461280 $Y=1036300
X1085 2864 1 2 2865 DELB $T=462520 981240 1 0 $X=462520 $Y=975820
X1086 2811 1 2 2848 DELB $T=463760 961080 0 0 $X=463760 $Y=960700
X1087 2901 1 2 2894 DELB $T=469960 900600 0 0 $X=469960 $Y=900220
X1088 2889 1 2 2917 DELB $T=473680 971160 0 0 $X=473680 $Y=970780
X1089 2929 1 2 2956 DELB $T=474920 1051800 0 0 $X=474920 $Y=1051420
X1090 2994 1 2 3010 DELB $T=486080 971160 1 0 $X=486080 $Y=965740
X1091 2965 1 2 2958 DELB $T=487940 940920 0 0 $X=487940 $Y=940540
X1092 3013 1 2 3050 DELB $T=494140 961080 1 0 $X=494140 $Y=955660
X1093 3021 1 2 3048 DELB $T=496000 930840 0 0 $X=496000 $Y=930460
X1094 3002 1 2 3076 DELB $T=499100 1061880 0 0 $X=499100 $Y=1061500
X1095 2986 1 2 3022 DELB $T=500340 1001400 1 0 $X=500340 $Y=995980
X1096 3057 1 2 3064 DELB $T=503440 1061880 1 0 $X=503440 $Y=1056460
X1097 3083 1 2 3046 DELB $T=504680 1021560 0 0 $X=504680 $Y=1021180
X1098 3073 1 2 3082 DELB $T=510260 951000 0 0 $X=510260 $Y=950620
X1099 3125 1 2 3128 DELB $T=510260 1061880 1 0 $X=510260 $Y=1056460
X1100 3091 1 2 3137 DELB $T=512740 1021560 0 0 $X=512740 $Y=1021180
X1101 3143 1 2 3145 DELB $T=514600 991320 1 0 $X=514600 $Y=985900
X1102 3153 1 2 3150 DELB $T=517080 1061880 1 0 $X=517080 $Y=1056460
X1103 3178 1 2 3179 DELB $T=520800 920760 1 0 $X=520800 $Y=915340
X1104 3188 1 2 3194 DELB $T=522660 951000 0 0 $X=522660 $Y=950620
X1105 3212 1 2 3211 DELB $T=527000 920760 1 0 $X=527000 $Y=915340
X1106 3207 1 2 3220 DELB $T=528240 1051800 0 0 $X=528240 $Y=1051420
X1107 3214 1 2 3243 DELB $T=533820 961080 1 0 $X=533820 $Y=955660
X1108 3318 1 2 3327 DELB $T=548080 920760 1 0 $X=548080 $Y=915340
X1109 3285 1 2 3362 DELB $T=554280 920760 1 0 $X=554280 $Y=915340
X1110 3308 1 2 3383 DELB $T=557380 1011480 0 0 $X=557380 $Y=1011100
X1111 3370 1 2 3367 DELB $T=561100 920760 0 0 $X=561100 $Y=920380
X1112 3423 1 2 3415 DELB $T=563580 1011480 1 0 $X=563580 $Y=1006060
X1113 3390 1 2 3432 DELB $T=565440 971160 0 0 $X=565440 $Y=970780
X1114 3365 1 2 3405 DELB $T=571020 940920 0 0 $X=571020 $Y=940540
X1115 3434 1 2 3422 DELB $T=571020 1011480 1 0 $X=571020 $Y=1006060
X1116 3468 1 2 3472 DELB $T=573500 981240 1 0 $X=573500 $Y=975820
X1117 3481 1 2 3460 DELB $T=575360 971160 1 0 $X=575360 $Y=965740
X1118 3478 1 2 3501 DELB $T=576600 940920 0 0 $X=576600 $Y=940540
X1119 3490 1 2 3515 DELB $T=580320 971160 0 0 $X=580320 $Y=970780
X1120 3529 1 2 3508 DELB $T=585280 930840 1 0 $X=585280 $Y=925420
X1121 3534 1 2 3533 DELB $T=585900 1021560 0 0 $X=585900 $Y=1021180
X1122 3520 1 2 3561 DELB $T=591480 930840 1 0 $X=591480 $Y=925420
X1123 3552 1 2 3555 DELB $T=592100 991320 0 0 $X=592100 $Y=990940
X1124 477 1 2 466 DELB $T=592720 900600 0 0 $X=592720 $Y=900220
X1125 3607 1 2 3634 DELB $T=603260 1001400 0 0 $X=603260 $Y=1001020
X1126 3619 1 2 3648 DELB $T=605120 1051800 1 0 $X=605120 $Y=1046380
X1127 3625 1 2 3630 DELB $T=606360 1071960 0 0 $X=606360 $Y=1071580
X1128 3641 1 2 3661 DELB $T=608220 1041720 0 0 $X=608220 $Y=1041340
X1129 3627 1 2 3651 DELB $T=611320 900600 0 0 $X=611320 $Y=900220
X1130 3660 1 2 3680 DELB $T=612560 1031640 0 0 $X=612560 $Y=1031260
X1131 3692 1 2 3719 DELB $T=617520 971160 0 0 $X=617520 $Y=970780
X1132 3670 1 2 3695 DELB $T=617520 1031640 1 0 $X=617520 $Y=1026220
X1133 3689 1 2 3712 DELB $T=620620 1082040 0 0 $X=620620 $Y=1081660
X1134 3738 1 2 3742 DELB $T=624340 1031640 1 0 $X=624340 $Y=1026220
X1135 3743 1 2 3769 DELB $T=629300 1061880 1 0 $X=629300 $Y=1056460
X1136 3771 1 2 3770 DELB $T=629300 1071960 0 0 $X=629300 $Y=1071580
X1137 3638 1 2 3729 DELB $T=631160 991320 0 0 $X=631160 $Y=990940
X1138 3764 1 2 3782 DELB $T=632400 1031640 1 0 $X=632400 $Y=1026220
X1139 3776 1 2 3797 DELB $T=634880 930840 0 0 $X=634880 $Y=930460
X1140 547 1 2 559 DELB $T=637360 1071960 0 0 $X=637360 $Y=1071580
X1141 3785 1 2 3780 DELB $T=638600 940920 0 0 $X=638600 $Y=940540
X1142 3791 1 2 3823 DELB $T=640460 1051800 1 0 $X=640460 $Y=1046380
X1143 3848 1 2 573 DELB $T=647280 900600 0 0 $X=647280 $Y=900220
X1144 3828 1 2 3847 DELB $T=647900 1031640 1 0 $X=647900 $Y=1026220
X1145 3829 1 2 3822 DELB $T=651000 1041720 1 0 $X=651000 $Y=1036300
X1146 571 1 2 584 DELB $T=653480 1082040 1 0 $X=653480 $Y=1076620
X1147 3873 1 2 3887 DELB $T=654720 951000 0 0 $X=654720 $Y=950620
X1148 3880 1 2 3915 DELB $T=656580 1041720 1 0 $X=656580 $Y=1036300
X1149 3906 1 2 3920 DELB $T=659680 1082040 1 0 $X=659680 $Y=1076620
X1150 3923 1 2 3931 DELB $T=668360 1051800 0 0 $X=668360 $Y=1051420
X1151 3919 1 2 3973 DELB $T=672700 1041720 0 0 $X=672700 $Y=1041340
X1152 3904 1 2 4016 DELB $T=673320 930840 1 0 $X=673320 $Y=925420
X1153 4009 1 2 4037 DELB $T=673940 1051800 0 0 $X=673940 $Y=1051420
X1154 4085 1 2 4118 DELB $T=686960 1031640 1 0 $X=686960 $Y=1026220
X1155 4048 1 2 4135 DELB $T=690680 920760 0 0 $X=690680 $Y=920380
X1156 4147 1 2 4179 DELB $T=697500 920760 1 0 $X=697500 $Y=915340
X1157 4125 1 2 4155 DELB $T=698120 1061880 0 0 $X=698120 $Y=1061500
X1158 4194 1 2 4218 DELB $T=704320 1021560 1 0 $X=704320 $Y=1016140
X1159 4203 1 2 4204 DELB $T=706180 930840 1 0 $X=706180 $Y=925420
X1160 4214 1 2 4251 DELB $T=710520 1082040 1 0 $X=710520 $Y=1076620
X1161 669 1 2 4261 DELB $T=717960 1071960 0 0 $X=717960 $Y=1071580
X1162 4309 1 2 4351 DELB $T=727260 930840 1 0 $X=727260 $Y=925420
X1163 4305 1 2 4342 DELB $T=729120 961080 0 0 $X=729120 $Y=960700
X1164 4334 1 2 4359 DELB $T=732220 1001400 0 0 $X=732220 $Y=1001020
X1165 4321 1 2 4371 DELB $T=734080 1082040 1 0 $X=734080 $Y=1076620
X1166 707 1 2 715 DELB $T=740900 910680 1 0 $X=740900 $Y=905260
X1167 4376 1 2 4389 DELB $T=744000 1051800 0 0 $X=744000 $Y=1051420
X1168 4386 1 2 4419 DELB $T=744620 1071960 0 0 $X=744620 $Y=1071580
X1169 4484 1 2 4462 DELB $T=759500 951000 0 0 $X=759500 $Y=950620
X1170 4492 1 2 4521 DELB $T=759500 1041720 1 0 $X=759500 $Y=1036300
X1171 4506 1 2 4529 DELB $T=761360 1041720 0 0 $X=761360 $Y=1041340
X1172 4517 1 2 4538 DELB $T=763220 940920 1 0 $X=763220 $Y=935500
X1173 4549 1 2 4583 DELB $T=769420 971160 1 0 $X=769420 $Y=965740
X1174 4581 1 2 4619 DELB $T=773760 1011480 0 0 $X=773760 $Y=1011100
X1175 4585 1 2 4584 DELB $T=773760 1051800 1 0 $X=773760 $Y=1046380
X1176 4610 1 2 4582 DELB $T=777480 940920 0 0 $X=777480 $Y=940540
X1177 4605 1 2 4651 DELB $T=778720 1082040 1 0 $X=778720 $Y=1076620
X1178 4625 1 2 4655 DELB $T=780580 981240 0 0 $X=780580 $Y=980860
X1179 4649 1 2 4681 DELB $T=784300 940920 0 0 $X=784300 $Y=940540
X1180 4648 1 2 4640 DELB $T=791120 910680 0 0 $X=791120 $Y=910300
X1181 4696 1 2 4730 DELB $T=791120 1041720 0 0 $X=791120 $Y=1041340
X1182 4617 1 2 4659 DELB $T=796700 991320 0 0 $X=796700 $Y=990940
X1183 4724 1 2 4731 DELB $T=798560 1071960 0 0 $X=798560 $Y=1071580
X1184 4805 1 2 4833 DELB $T=806620 1071960 0 0 $X=806620 $Y=1071580
X1185 4818 1 2 4849 DELB $T=807860 951000 1 0 $X=807860 $Y=945580
X1186 4839 1 2 4840 DELB $T=814680 991320 1 0 $X=814680 $Y=985900
X1187 4879 1 2 4906 DELB $T=817160 910680 1 0 $X=817160 $Y=905260
X1188 4845 1 2 4855 DELB $T=819020 961080 0 0 $X=819020 $Y=960700
X1189 4860 1 2 4895 DELB $T=819640 1082040 0 0 $X=819640 $Y=1081660
X1190 4901 1 2 4900 DELB $T=821500 940920 0 0 $X=821500 $Y=940540
X1191 4946 1 2 4949 DELB $T=831420 971160 0 0 $X=831420 $Y=970780
X1192 4960 1 2 4986 DELB $T=833900 910680 1 0 $X=833900 $Y=905260
X1193 4873 1 2 4945 DELB $T=835140 1051800 0 0 $X=835140 $Y=1051420
X1194 4974 1 2 4980 DELB $T=836380 930840 0 0 $X=836380 $Y=930460
X1195 5003 1 2 4989 DELB $T=841340 910680 0 0 $X=841340 $Y=910300
X1196 5001 1 2 5043 DELB $T=847540 951000 1 0 $X=847540 $Y=945580
X1197 5045 1 2 5044 DELB $T=847540 1021560 1 0 $X=847540 $Y=1016140
X1198 5048 1 2 5049 DELB $T=848160 910680 0 0 $X=848160 $Y=910300
X1199 5051 1 2 5071 DELB $T=848160 1001400 1 0 $X=848160 $Y=995980
X1200 5068 1 2 5030 DELB $T=851260 1051800 0 0 $X=851260 $Y=1051420
X1201 5069 1 2 5080 DELB $T=854360 1021560 1 0 $X=854360 $Y=1016140
X1202 5100 1 2 5087 DELB $T=857460 971160 1 0 $X=857460 $Y=965740
X1203 5094 1 2 5118 DELB $T=860560 1021560 1 0 $X=860560 $Y=1016140
X1204 5128 1 2 5122 DELB $T=862420 971160 0 0 $X=862420 $Y=970780
X1205 5185 1 2 5150 DELB $T=876680 1001400 0 0 $X=876680 $Y=1001020
X1206 5222 1 2 5237 DELB $T=879780 930840 0 0 $X=879780 $Y=930460
X1207 5281 1 2 5273 DELB $T=885980 961080 1 0 $X=885980 $Y=955660
X1208 5276 1 2 5291 DELB $T=891560 1082040 0 0 $X=891560 $Y=1081660
X1209 5130 1 2 5121 DELB $T=892180 971160 0 0 $X=892180 $Y=970780
X1210 5327 1 2 5334 DELB $T=894040 1011480 0 0 $X=894040 $Y=1011100
X1211 5244 1 2 5289 DELB $T=894660 1061880 0 0 $X=894660 $Y=1061500
X1212 5351 1 2 5349 DELB $T=897140 1051800 0 0 $X=897140 $Y=1051420
X1213 5187 1 2 5301 DELB $T=899620 1082040 0 0 $X=899620 $Y=1081660
X1214 5221 1 2 5190 DELB $T=901480 951000 0 0 $X=901480 $Y=950620
X1215 5302 1 2 5326 DELB $T=902720 910680 0 0 $X=902720 $Y=910300
X1216 5427 1 2 5445 DELB $T=919460 1051800 0 0 $X=919460 $Y=1051420
X1217 976 1 2 988 DELB $T=919460 1082040 0 0 $X=919460 $Y=1081660
X1218 5423 1 2 5441 DELB $T=923180 1001400 1 0 $X=923180 $Y=995980
X1219 5443 1 2 5444 DELB $T=923180 1051800 1 0 $X=923180 $Y=1046380
X1220 5484 1 2 5516 DELB $T=925040 900600 0 0 $X=925040 $Y=900220
X1221 5104 1 2 5133 DELB $T=925040 961080 1 0 $X=925040 $Y=955660
X1222 5515 1 2 5514 DELB $T=930620 1051800 1 0 $X=930620 $Y=1046380
X1223 5561 1 2 5596 DELB $T=938680 1021560 1 0 $X=938680 $Y=1016140
X1224 1017 1 2 1024 DELB $T=939920 900600 0 0 $X=939920 $Y=900220
X1225 5544 1 2 5580 DELB $T=940540 920760 1 0 $X=940540 $Y=915340
X1226 1015 1 2 5584 DELB $T=941160 1082040 1 0 $X=941160 $Y=1076620
X1227 5522 1 2 5555 DELB $T=942400 1031640 0 0 $X=942400 $Y=1031260
X1228 5615 1 2 5653 DELB $T=947360 971160 0 0 $X=947360 $Y=970780
X1229 5641 1 2 5633 DELB $T=951700 1031640 0 0 $X=951700 $Y=1031260
X1230 5590 1 2 5605 DELB $T=954180 930840 0 0 $X=954180 $Y=930460
X1231 5677 1 2 5676 DELB $T=956660 1082040 1 0 $X=956660 $Y=1076620
X1232 5672 1 2 5667 DELB $T=958520 961080 1 0 $X=958520 $Y=955660
X1233 5658 1 2 5692 DELB $T=959140 1031640 0 0 $X=959140 $Y=1031260
X1234 5629 1 2 5607 DELB $T=959760 991320 1 0 $X=959760 $Y=985900
X1235 5691 1 2 5727 DELB $T=965340 961080 1 0 $X=965340 $Y=955660
X1236 5724 1 2 5728 DELB $T=965340 991320 1 0 $X=965340 $Y=985900
X1237 5776 1 2 5795 DELB $T=981460 991320 0 0 $X=981460 $Y=990940
X1238 5778 1 2 5749 DELB $T=984560 961080 1 0 $X=984560 $Y=955660
X1239 1075 1 2 5843 DELB $T=987040 1082040 0 0 $X=987040 $Y=1081660
X1240 5824 1 2 5827 DELB $T=987660 900600 0 0 $X=987660 $Y=900220
X1241 5842 1 2 5864 DELB $T=991380 1071960 0 0 $X=991380 $Y=1071580
X1242 5885 1 2 5917 DELB $T=1000680 910680 0 0 $X=1000680 $Y=910300
X1243 5889 1 2 5871 DELB $T=1005640 910680 1 0 $X=1005640 $Y=905260
X1244 5932 1 2 5909 DELB $T=1005640 1021560 1 0 $X=1005640 $Y=1016140
X1245 5868 1 2 5888 DELB $T=1008120 1071960 0 0 $X=1008120 $Y=1071580
X1246 5957 1 2 5992 DELB $T=1011220 951000 0 0 $X=1011220 $Y=950620
X1247 5987 1 2 5988 DELB $T=1015560 910680 1 0 $X=1015560 $Y=905260
X1248 5965 1 2 6005 DELB $T=1018660 1041720 0 0 $X=1018660 $Y=1041340
X1249 5985 1 2 5999 DELB $T=1023000 1001400 1 0 $X=1023000 $Y=995980
X1250 6022 1 2 6059 DELB $T=1029200 1082040 1 0 $X=1029200 $Y=1076620
X1251 6074 1 2 6100 DELB $T=1032300 940920 1 0 $X=1032300 $Y=935500
X1252 6023 1 2 6086 DELB $T=1034160 1001400 1 0 $X=1034160 $Y=995980
X1253 6015 1 2 6051 DELB $T=1035400 1041720 0 0 $X=1035400 $Y=1041340
X1254 5982 1 2 5949 DELB $T=1037880 910680 0 0 $X=1037880 $Y=910300
X1255 6025 1 2 6058 DELB $T=1039120 951000 0 0 $X=1039120 $Y=950620
X1256 6124 1 2 6133 DELB $T=1042220 1031640 0 0 $X=1042220 $Y=1031260
X1257 6036 1 2 6061 DELB $T=1048420 1031640 0 0 $X=1048420 $Y=1031260
X1258 6165 1 2 6189 DELB $T=1050900 920760 0 0 $X=1050900 $Y=920380
X1259 6134 1 2 6164 DELB $T=1054000 1061880 0 0 $X=1054000 $Y=1061500
X1260 1189 1 2 1199 DELB $T=1055860 1082040 0 0 $X=1055860 $Y=1081660
X1261 6138 1 2 6136 DELB $T=1056480 1011480 1 0 $X=1056480 $Y=1006060
X1262 6225 1 2 6238 DELB $T=1063300 1011480 1 0 $X=1063300 $Y=1006060
X1263 6243 1 2 6269 DELB $T=1064540 1021560 1 0 $X=1064540 $Y=1016140
X1264 6209 1 2 6239 DELB $T=1065160 1041720 1 0 $X=1065160 $Y=1036300
X1265 6035 1 2 6089 DELB $T=1073840 1001400 0 0 $X=1073840 $Y=1001020
X1266 6284 1 2 6279 DELB $T=1076320 1031640 0 0 $X=1076320 $Y=1031260
X1267 1222 1 2 1229 DELB $T=1079420 900600 0 0 $X=1079420 $Y=900220
X1268 6322 1 2 6329 DELB $T=1081900 1061880 1 0 $X=1081900 $Y=1056460
X1269 1242 1 2 1249 DELB $T=1093680 910680 1 0 $X=1093680 $Y=905260
X1270 6373 1 2 6368 DELB $T=1096780 1031640 1 0 $X=1096780 $Y=1026220
X1271 6413 1 2 6432 DELB $T=1098640 930840 0 0 $X=1098640 $Y=930460
X1272 6414 1 2 6449 DELB $T=1102360 991320 0 0 $X=1102360 $Y=990940
X1273 6411 1 2 6437 DELB $T=1104220 1031640 1 0 $X=1104220 $Y=1026220
X1274 6446 1 2 6473 DELB $T=1106080 1051800 0 0 $X=1106080 $Y=1051420
X1275 6453 1 2 6479 DELB $T=1109180 991320 0 0 $X=1109180 $Y=990940
X1276 6463 1 2 6470 DELB $T=1110420 1071960 0 0 $X=1110420 $Y=1071580
X1277 6430 1 2 6475 DELB $T=1111040 930840 0 0 $X=1111040 $Y=930460
X1278 6461 1 2 6502 DELB $T=1111040 951000 0 0 $X=1111040 $Y=950620
X1279 1278 1 2 6466 DELB $T=1113520 1082040 0 0 $X=1113520 $Y=1081660
X1280 6439 1 2 6478 DELB $T=1116000 951000 1 0 $X=1116000 $Y=945580
X1281 6505 1 2 6520 DELB $T=1117860 930840 0 0 $X=1117860 $Y=930460
X1282 6433 1 2 6474 DELB $T=1120340 900600 0 0 $X=1120340 $Y=900220
X1283 6506 1 2 6519 DELB $T=1121580 1001400 0 0 $X=1121580 $Y=1001020
X1284 6448 1 2 6483 DELB $T=1123440 1082040 0 0 $X=1123440 $Y=1081660
X1285 6509 1 2 6525 DELB $T=1124680 951000 1 0 $X=1124680 $Y=945580
X1286 1350 1 2 1345 DELA $T=230020 1011480 0 0 $X=230020 $Y=1011100
X1287 1397 1 2 1405 DELA $T=234360 1021560 1 0 $X=234360 $Y=1016140
X1288 1446 1 2 1472 DELA $T=241180 1011480 1 0 $X=241180 $Y=1006060
X1289 1386 1 2 1339 DELA $T=249240 991320 0 0 $X=249240 $Y=990940
X1290 1643 1 2 1638 DELA $T=272180 1021560 0 0 $X=272180 $Y=1021180
X1291 1724 1 2 1804 DELA $T=294500 991320 1 0 $X=294500 $Y=985900
X1292 1514 1 2 1767 DELA $T=296980 1021560 1 0 $X=296980 $Y=1016140
X1293 74 1 2 1877 DELA $T=299460 991320 1 0 $X=299460 $Y=985900
X1294 1950 1 2 1948 DELA $T=314960 981240 0 0 $X=314960 $Y=980860
X1295 1984 1 2 1978 DELA $T=322400 1011480 1 0 $X=322400 $Y=1006060
X1296 126 1 2 2053 DELA $T=327980 1011480 1 0 $X=327980 $Y=1006060
X1297 134 1 2 2090 DELA $T=332940 1011480 1 0 $X=332940 $Y=1006060
X1298 132 1 2 2044 DELA $T=332940 1031640 0 0 $X=332940 $Y=1031260
X1299 137 1 2 2093 DELA $T=337900 1011480 1 0 $X=337900 $Y=1006060
X1300 2096 1 2 2128 DELA $T=338520 981240 1 0 $X=338520 $Y=975820
X1301 151 1 2 2160 DELA $T=343480 1011480 1 0 $X=343480 $Y=1006060
X1302 2123 1 2 2165 DELA $T=344100 971160 1 0 $X=344100 $Y=965740
X1303 2189 1 2 2217 DELA $T=352160 981240 1 0 $X=352160 $Y=975820
X1304 2219 1 2 2241 DELA $T=356500 1031640 0 0 $X=356500 $Y=1031260
X1305 2231 1 2 2250 DELA $T=358980 981240 0 0 $X=358980 $Y=980860
X1306 1669 1 2 2251 DELA $T=363320 1071960 1 0 $X=363320 $Y=1066540
X1307 2256 1 2 2287 DELA $T=363940 981240 0 0 $X=363940 $Y=980860
X1308 2261 1 2 2295 DELA $T=365180 951000 1 0 $X=365180 $Y=945580
X1309 2272 1 2 2304 DELA $T=366420 971160 0 0 $X=366420 $Y=970780
X1310 2365 1 2 2392 DELA $T=379440 930840 0 0 $X=379440 $Y=930460
X1311 2382 1 2 2408 DELA $T=382540 981240 1 0 $X=382540 $Y=975820
X1312 2410 1 2 2437 DELA $T=386880 940920 1 0 $X=386880 $Y=935500
X1313 2413 1 2 2444 DELA $T=387500 981240 1 0 $X=387500 $Y=975820
X1314 2452 1 2 2459 DELA $T=392460 981240 1 0 $X=392460 $Y=975820
X1315 2458 1 2 2480 DELA $T=393700 940920 1 0 $X=393700 $Y=935500
X1316 2509 1 2 2545 DELA $T=403620 951000 0 0 $X=403620 $Y=950620
X1317 224 1 2 228 DELA $T=404860 900600 0 0 $X=404860 $Y=900220
X1318 2532 1 2 2558 DELA $T=406100 930840 1 0 $X=406100 $Y=925420
X1319 229 1 2 233 DELA $T=409820 900600 0 0 $X=409820 $Y=900220
X1320 2584 1 2 2618 DELA $T=414780 920760 1 0 $X=414780 $Y=915340
X1321 2551 1 2 2606 DELA $T=417260 981240 0 0 $X=417260 $Y=980860
X1322 2612 1 2 2613 DELA $T=419120 951000 1 0 $X=419120 $Y=945580
X1323 2639 1 2 2656 DELA $T=425320 981240 0 0 $X=425320 $Y=980860
X1324 2662 1 2 2708 DELA $T=430900 951000 0 0 $X=430900 $Y=950620
X1325 2729 1 2 2695 DELA $T=441440 971160 1 0 $X=441440 $Y=965740
X1326 2830 1 2 2831 DELA $T=456320 981240 1 0 $X=456320 $Y=975820
X1327 2916 1 2 2915 DELA $T=472440 961080 0 0 $X=472440 $Y=960700
X1328 2911 1 2 2890 DELA $T=478640 971160 1 0 $X=478640 $Y=965740
X1329 2933 1 2 2943 DELA $T=510880 1001400 0 0 $X=510880 $Y=1001020
X1330 3156 1 2 3142 DELA $T=517700 951000 0 0 $X=517700 $Y=950620
X1331 329 1 2 3043 DELA $T=527620 940920 1 0 $X=527620 $Y=935500
X1332 3299 1 2 3300 DELA $T=543120 930840 1 0 $X=543120 $Y=925420
X1333 3599 1 2 3618 DELA $T=600780 961080 0 0 $X=600780 $Y=960700
X1334 3639 1 2 3659 DELA $T=608220 1001400 0 0 $X=608220 $Y=1001020
X1335 3694 1 2 3693 DELA $T=617520 1001400 0 0 $X=617520 $Y=1001020
X1336 3808 1 2 3827 DELA $T=638600 991320 0 0 $X=638600 $Y=990940
X1337 3790 1 2 3831 DELA $T=639220 1021560 0 0 $X=639220 $Y=1021180
X1338 3851 1 2 3876 DELA $T=647900 991320 1 0 $X=647900 $Y=985900
X1339 4095 1 2 4133 DELA $T=694400 981240 0 0 $X=694400 $Y=980860
X1340 4266 1 2 4298 DELA $T=719820 991320 0 0 $X=719820 $Y=990940
X1341 4320 1 2 4354 DELA $T=727260 1001400 0 0 $X=727260 $Y=1001020
X1342 4235 1 2 4200 DELA $T=734080 961080 0 0 $X=734080 $Y=960700
X1343 4510 1 2 4530 DELA $T=761980 1011480 0 0 $X=761980 $Y=1011100
X1344 4554 1 2 4587 DELA $T=770040 930840 0 0 $X=770040 $Y=930460
X1345 4793 1 2 4798 DELA $T=822740 1031640 0 0 $X=822740 $Y=1031260
X1346 5088 1 2 5119 DELA $T=856840 1051800 0 0 $X=856840 $Y=1051420
X1347 5155 1 2 5156 DELA $T=866760 1021560 1 0 $X=866760 $Y=1016140
X1348 5377 1 2 5384 DELA $T=903960 1061880 1 0 $X=903960 $Y=1056460
X1349 5325 1 2 5347 DELA $T=905820 1031640 1 0 $X=905820 $Y=1026220
X1350 5393 1 2 5408 DELA $T=905820 1082040 0 0 $X=905820 $Y=1081660
X1351 5556 1 2 5587 DELA $T=937440 1051800 0 0 $X=937440 $Y=1051420
X1352 5647 1 2 5674 DELA $T=951080 1031640 1 0 $X=951080 $Y=1026220
X1353 5819 1 2 5835 DELA $T=986420 920760 0 0 $X=986420 $Y=920380
X1354 5823 1 2 5839 DELA $T=987040 971160 1 0 $X=987040 $Y=965740
X1355 5836 1 2 5862 DELA $T=990760 981240 0 0 $X=990760 $Y=980860
X1356 5929 1 2 5931 DELA $T=1005640 951000 0 0 $X=1005640 $Y=950620
X1357 5960 1 2 5997 DELA $T=1016800 991320 0 0 $X=1016800 $Y=990940
X1358 5886 1 2 5946 DELA $T=1019900 940920 1 0 $X=1019900 $Y=935500
X1359 6040 1 2 6057 DELA $T=1027340 940920 1 0 $X=1027340 $Y=935500
X1360 6139 1 2 6140 DELA $T=1044700 920760 0 0 $X=1044700 $Y=920380
X1361 6122 1 2 6170 DELA $T=1051520 1011480 1 0 $X=1051520 $Y=1006060
X1362 6135 1 2 1196 DELA $T=1055240 920760 1 0 $X=1055240 $Y=915340
X1363 6213 1 2 6235 DELA $T=1067020 920760 0 0 $X=1067020 $Y=920380
X1364 6405 1 2 6420 DELA $T=1097400 991320 0 0 $X=1097400 $Y=990940
X1365 6343 1 2 6361 DELA $T=1102360 951000 0 0 $X=1102360 $Y=950620
X1366 1281 1 2 1284 DELA $T=1118480 1082040 0 0 $X=1118480 $Y=1081660
X1367 6452 1 2 6467 DELA $T=1119100 961080 0 0 $X=1119100 $Y=960700
X1368 6376 1 2 6375 DELA $T=1124060 961080 0 0 $X=1124060 $Y=960700
X1369 1308 4 1358 2 1 1350 QDFFRBN $T=220720 1001400 0 0 $X=220720 $Y=1001020
X1370 1316 4 1358 2 1 1338 QDFFRBN $T=221340 981240 0 0 $X=221340 $Y=980860
X1371 1317 4 1358 2 1 1386 QDFFRBN $T=221340 991320 0 0 $X=221340 $Y=990940
X1372 1395 4 1358 2 1 1397 QDFFRBN $T=233740 1001400 0 0 $X=233740 $Y=1001020
X1373 1442 4 1358 2 1 1402 QDFFRBN $T=246760 981240 1 180 $X=234980 $Y=980860
X1374 1477 4 1358 2 1 1447 QDFFRBN $T=253580 991320 0 180 $X=241800 $Y=985900
X1375 1537 4 1451 2 1 1446 QDFFRBN $T=259160 1001400 1 180 $X=247380 $Y=1001020
X1376 1533 4 1451 2 1 1608 QDFFRBN $T=253580 1011480 1 0 $X=253580 $Y=1006060
X1377 1582 4 1451 2 1 1630 QDFFRBN $T=261020 1001400 0 0 $X=261020 $Y=1001020
X1378 1626 4 1451 2 1 1644 QDFFRBN $T=267840 1011480 1 0 $X=267840 $Y=1006060
X1379 1745 4 1451 2 1 1554 QDFFRBN $T=287060 1001400 1 180 $X=275280 $Y=1001020
X1380 1791 4 1716 2 1 1724 QDFFRBN $T=293880 1011480 0 180 $X=282100 $Y=1006060
X1381 1787 4 1716 2 1 1514 QDFFRBN $T=294500 1011480 1 180 $X=282720 $Y=1011100
X1382 1793 4 75 2 1 1870 QDFFRBN $T=292020 1082040 0 0 $X=292020 $Y=1081660
X1383 1888 4 1716 2 1 1796 QDFFRBN $T=306900 1001400 1 180 $X=295120 $Y=1001020
X1384 1810 4 1716 2 1 1541 QDFFRBN $T=297600 1011480 0 0 $X=297600 $Y=1011100
X1385 1836 4 1716 2 1 1912 QDFFRBN $T=297600 1021560 0 0 $X=297600 $Y=1021180
X1386 1916 4 75 2 1 1950 QDFFRBN $T=309380 1011480 1 0 $X=309380 $Y=1006060
X1387 1924 4 1910 2 1 1989 QDFFRBN $T=311860 991320 1 0 $X=311860 $Y=985900
X1388 1932 4 1910 2 1 1997 QDFFRBN $T=312480 991320 0 0 $X=312480 $Y=990940
X1389 1933 4 1976 2 1 1988 QDFFRBN $T=312480 1021560 0 0 $X=312480 $Y=1021180
X1390 1927 4 1910 2 1 1944 QDFFRBN $T=313720 981240 1 0 $X=313720 $Y=975820
X1391 1966 4 1910 2 1 1984 QDFFRBN $T=318060 1001400 0 0 $X=318060 $Y=1001020
X1392 1990 4 1976 2 1 2024 QDFFRBN $T=323020 1011480 0 0 $X=323020 $Y=1011100
X1393 2070 4 1976 2 1 132 QDFFRBN $T=343480 1021560 1 180 $X=331700 $Y=1021180
X1394 2056 4 1976 2 1 126 QDFFRBN $T=332320 1001400 0 0 $X=332320 $Y=1001020
X1395 2084 4 1976 2 1 137 QDFFRBN $T=347820 1021560 0 180 $X=336040 $Y=1016140
X1396 2118 4 2184 2 1 2175 QDFFRBN $T=343480 1071960 0 0 $X=343480 $Y=1071580
X1397 2140 4 2184 2 1 2109 QDFFRBN $T=344100 1061880 0 0 $X=344100 $Y=1061500
X1398 2145 4 2184 2 1 2146 QDFFRBN $T=345960 1061880 1 0 $X=345960 $Y=1056460
X1399 2164 4 2184 2 1 2163 QDFFRBN $T=349680 1051800 0 0 $X=349680 $Y=1051420
X1400 175 4 168 2 1 161 QDFFRBN $T=362080 1082040 1 180 $X=350300 $Y=1081660
X1401 2180 4 2233 2 1 2210 QDFFRBN $T=350920 1011480 0 0 $X=350920 $Y=1011100
X1402 2186 4 1976 2 1 2096 QDFFRBN $T=351540 1001400 1 0 $X=351540 $Y=995980
X1403 2216 4 2258 2 1 2292 QDFFRBN $T=355880 1071960 0 0 $X=355880 $Y=1071580
X1404 2208 4 2184 2 1 2220 QDFFRBN $T=357120 1041720 0 0 $X=357120 $Y=1041340
X1405 2227 4 2275 2 1 2260 QDFFRBN $T=358360 1061880 0 0 $X=358360 $Y=1061500
X1406 2254 4 2233 2 1 134 QDFFRBN $T=363320 1021560 1 0 $X=363320 $Y=1016140
X1407 2277 185 2334 2 1 2356 QDFFRBN $T=366420 1051800 0 0 $X=366420 $Y=1051420
X1408 2278 185 2275 2 1 2355 QDFFRBN $T=366420 1061880 1 0 $X=366420 $Y=1056460
X1409 2285 185 2258 2 1 2330 QDFFRBN $T=367660 1082040 1 0 $X=367660 $Y=1076620
X1410 2302 185 2275 2 1 2374 QDFFRBN $T=370140 1041720 0 0 $X=370140 $Y=1041340
X1411 2303 185 2258 2 1 2381 QDFFRBN $T=370140 1071960 1 0 $X=370140 $Y=1066540
X1412 2336 185 2380 2 1 2390 QDFFRBN $T=374480 1021560 0 0 $X=374480 $Y=1021180
X1413 2034 185 2394 2 1 2317 QDFFRBN $T=375720 991320 0 0 $X=375720 $Y=990940
X1414 2347 185 2233 2 1 151 QDFFRBN $T=389360 1011480 1 180 $X=377580 $Y=1011100
X1415 2362 185 2379 2 1 2243 QDFFRBN $T=378200 1021560 1 0 $X=378200 $Y=1016140
X1416 2424 185 2275 2 1 2329 QDFFRBN $T=391220 1061880 0 180 $X=379440 $Y=1056460
X1417 2422 185 2380 2 1 2452 QDFFRBN $T=389360 991320 0 0 $X=389360 $Y=990940
X1418 2423 185 2380 2 1 2383 QDFFRBN $T=389360 1001400 1 0 $X=389360 $Y=995980
X1419 2441 185 2379 2 1 2520 QDFFRBN $T=390600 1011480 1 0 $X=390600 $Y=1006060
X1420 2443 185 2334 2 1 2457 QDFFRBN $T=391220 1051800 1 0 $X=391220 $Y=1046380
X1421 2494 185 2334 2 1 2440 QDFFRBN $T=403000 1061880 1 180 $X=391220 $Y=1061500
X1422 2453 185 2492 2 1 2461 QDFFRBN $T=392460 1011480 0 0 $X=392460 $Y=1011100
X1423 2460 185 2334 2 1 2313 QDFFRBN $T=393700 1061880 1 0 $X=393700 $Y=1056460
X1424 2511 185 2379 2 1 2300 QDFFRBN $T=407960 1031640 1 180 $X=396180 $Y=1031260
X1425 2543 185 2394 2 1 2458 QDFFRBN $T=409200 971160 0 180 $X=397420 $Y=965740
X1426 2481 185 2394 2 1 2290 QDFFRBN $T=398040 991320 1 0 $X=398040 $Y=985900
X1427 2514 185 2492 2 1 2348 QDFFRBN $T=412920 1021560 0 180 $X=401140 $Y=1016140
X1428 2594 185 2394 2 1 2498 QDFFRBN $T=414160 971160 1 180 $X=402380 $Y=970780
X1429 2508 185 2394 2 1 2501 QDFFRBN $T=403000 1001400 1 0 $X=403000 $Y=995980
X1430 2599 185 2492 2 1 2534 QDFFRBN $T=417880 1021560 1 180 $X=406100 $Y=1021180
X1431 2608 185 2334 2 1 2541 QDFFRBN $T=419120 1061880 0 180 $X=407340 $Y=1056460
X1432 2617 185 2570 2 1 2551 QDFFRBN $T=420980 991320 1 180 $X=409200 $Y=990940
X1433 2555 185 2492 2 1 2526 QDFFRBN $T=409200 1031640 0 0 $X=409200 $Y=1031260
X1434 2622 185 2492 2 1 2516 QDFFRBN $T=421600 1011480 0 180 $X=409820 $Y=1006060
X1435 2565 185 2570 2 1 2638 QDFFRBN $T=411060 971160 1 0 $X=411060 $Y=965740
X1436 2567 185 2614 2 1 2493 QDFFRBN $T=411680 1041720 0 0 $X=411680 $Y=1041340
X1437 2641 185 2492 2 1 2611 QDFFRBN $T=430280 1011480 1 180 $X=418500 $Y=1011100
X1438 2623 185 2614 2 1 2658 QDFFRBN $T=419740 1041720 1 0 $X=419740 $Y=1036300
X1439 2628 2637 2651 2 1 2612 QDFFRBN $T=420360 961080 0 0 $X=420360 $Y=960700
X1440 2629 185 2644 2 1 2694 QDFFRBN $T=420360 1021560 0 0 $X=420360 $Y=1021180
X1441 2630 185 2614 2 1 2668 QDFFRBN $T=420360 1051800 0 0 $X=420360 $Y=1051420
X1442 2635 185 236 2 1 2647 QDFFRBN $T=420980 1082040 1 0 $X=420980 $Y=1076620
X1443 2700 252 236 2 1 242 QDFFRBN $T=434620 1082040 1 180 $X=422840 $Y=1081660
X1444 2648 185 2570 2 1 2729 QDFFRBN $T=423460 991320 0 0 $X=423460 $Y=990940
X1445 2659 2637 2570 2 1 2704 QDFFRBN $T=425320 971160 1 0 $X=425320 $Y=965740
X1446 2720 2637 2651 2 1 2662 QDFFRBN $T=437720 961080 0 180 $X=425940 $Y=955660
X1447 2725 2637 2570 2 1 2382 QDFFRBN $T=442060 991320 0 180 $X=430280 $Y=985900
X1448 2690 253 2734 2 1 2703 QDFFRBN $T=430900 940920 1 0 $X=430900 $Y=935500
X1449 2691 185 2644 2 1 2757 QDFFRBN $T=430900 1001400 0 0 $X=430900 $Y=1001020
X1450 2697 2637 2651 2 1 2743 QDFFRBN $T=432140 971160 0 0 $X=432140 $Y=970780
X1451 2699 185 262 2 1 2772 QDFFRBN $T=432760 1061880 0 0 $X=432760 $Y=1061500
X1452 2706 253 263 2 1 2726 QDFFRBN $T=434000 910680 0 0 $X=434000 $Y=910300
X1453 2764 2637 2644 2 1 2705 QDFFRBN $T=445780 1021560 1 180 $X=434000 $Y=1021180
X1454 2707 185 262 2 1 2667 QDFFRBN $T=434000 1051800 0 0 $X=434000 $Y=1051420
X1455 256 253 263 2 1 2717 QDFFRBN $T=434620 900600 0 0 $X=434620 $Y=900220
X1456 2715 253 263 2 1 2687 QDFFRBN $T=435240 920760 1 0 $X=435240 $Y=915340
X1457 2719 253 2753 2 1 2410 QDFFRBN $T=435860 930840 0 0 $X=435860 $Y=930460
X1458 2760 2637 2644 2 1 2689 QDFFRBN $T=448260 1011480 0 180 $X=436480 $Y=1006060
X1459 2739 2637 2734 2 1 2722 QDFFRBN $T=439580 961080 0 0 $X=439580 $Y=960700
X1460 2746 253 2753 2 1 275 QDFFRBN $T=441440 930840 1 0 $X=441440 $Y=925420
X1461 2756 2637 2734 2 1 2776 QDFFRBN $T=443920 991320 1 0 $X=443920 $Y=985900
X1462 2758 252 2806 2 1 271 QDFFRBN $T=443920 1082040 1 0 $X=443920 $Y=1076620
X1463 2755 252 2806 2 1 2589 QDFFRBN $T=443920 1082040 0 0 $X=443920 $Y=1081660
X1464 2769 253 263 2 1 281 QDFFRBN $T=445780 910680 1 0 $X=445780 $Y=905260
X1465 2773 253 2753 2 1 2817 QDFFRBN $T=446400 940920 1 0 $X=446400 $Y=935500
X1466 2787 2637 2828 2 1 2809 QDFFRBN $T=447640 1021560 1 0 $X=447640 $Y=1016140
X1467 2788 252 262 2 1 2834 QDFFRBN $T=447640 1041720 0 0 $X=447640 $Y=1041340
X1468 2804 252 262 2 1 2709 QDFFRBN $T=459420 1051800 1 180 $X=447640 $Y=1051420
X1469 2791 253 279 2 1 2853 QDFFRBN $T=448260 910680 0 0 $X=448260 $Y=910300
X1470 2794 252 2806 2 1 2740 QDFFRBN $T=448880 1071960 1 0 $X=448880 $Y=1066540
X1471 2766 2637 2828 2 1 2274 QDFFRBN $T=451360 1011480 0 0 $X=451360 $Y=1011100
X1472 2814 2637 2825 2 1 2833 QDFFRBN $T=453220 971160 0 0 $X=453220 $Y=970780
X1473 2816 253 2875 2 1 2742 QDFFRBN $T=456320 930840 1 0 $X=456320 $Y=925420
X1474 2841 252 2806 2 1 2869 QDFFRBN $T=457560 1082040 1 0 $X=457560 $Y=1076620
X1475 2868 2637 2825 2 1 2811 QDFFRBN $T=470580 971160 0 180 $X=458800 $Y=965740
X1476 2852 253 279 2 1 2901 QDFFRBN $T=460040 910680 1 0 $X=460040 $Y=905260
X1477 2850 2637 2828 2 1 2864 QDFFRBN $T=460040 991320 0 0 $X=460040 $Y=990940
X1478 2863 2637 2875 2 1 2797 QDFFRBN $T=473060 951000 1 180 $X=461280 $Y=950620
X1479 2893 252 2876 2 1 2798 QDFFRBN $T=473060 1051800 1 180 $X=461280 $Y=1051420
X1480 2861 252 2876 2 1 300 QDFFRBN $T=461900 1041720 0 0 $X=461900 $Y=1041340
X1481 2870 2637 2828 2 1 2907 QDFFRBN $T=463140 1021560 0 0 $X=463140 $Y=1021180
X1482 2821 252 2876 2 1 2843 QDFFRBN $T=474920 1051800 0 180 $X=463140 $Y=1046380
X1483 2922 2637 2875 2 1 2438 QDFFRBN $T=475540 961080 0 180 $X=463760 $Y=955660
X1484 2897 252 2806 2 1 2872 QDFFRBN $T=475540 1061880 1 180 $X=463760 $Y=1061500
X1485 2883 253 2753 2 1 2916 QDFFRBN $T=465620 940920 1 0 $X=465620 $Y=935500
X1486 2885 2637 2887 2 1 2911 QDFFRBN $T=466240 1011480 0 0 $X=466240 $Y=1011100
X1487 2935 2637 2825 2 1 2889 QDFFRBN $T=479880 981240 0 180 $X=468100 $Y=975820
X1488 2899 2637 2941 2 1 2962 QDFFRBN $T=469340 951000 1 0 $X=469340 $Y=945580
X1489 2910 2637 2828 2 1 2949 QDFFRBN $T=470580 1001400 1 0 $X=470580 $Y=995980
X1490 2914 253 2951 2 1 2975 QDFFRBN $T=471200 930840 1 0 $X=471200 $Y=925420
X1491 2909 252 2944 2 1 2920 QDFFRBN $T=471200 1082040 1 0 $X=471200 $Y=1076620
X1492 2923 2637 2887 2 1 2987 QDFFRBN $T=473680 1011480 1 0 $X=473680 $Y=1006060
X1493 2964 253 2951 2 1 2660 QDFFRBN $T=487940 910680 0 180 $X=476160 $Y=905260
X1494 2952 252 2876 2 1 301 QDFFRBN $T=487940 1041720 1 180 $X=476160 $Y=1041340
X1495 2960 2637 2887 2 1 2933 QDFFRBN $T=488560 1021560 1 180 $X=476780 $Y=1021180
X1496 2946 2637 2941 2 1 2548 QDFFRBN $T=477400 961080 0 0 $X=477400 $Y=960700
X1497 2953 252 2944 2 1 2973 QDFFRBN $T=478640 1061880 0 0 $X=478640 $Y=1061500
X1498 323 253 2951 2 1 308 QDFFRBN $T=491660 900600 1 180 $X=479880 $Y=900220
X1499 3014 2637 2955 2 1 2959 QDFFRBN $T=491660 981240 1 180 $X=479880 $Y=980860
X1500 2998 252 2950 2 1 2929 QDFFRBN $T=491660 1051800 0 180 $X=479880 $Y=1046380
X1501 2966 2637 2941 2 1 2222 QDFFRBN $T=480500 951000 0 0 $X=480500 $Y=950620
X1502 3015 2637 2955 2 1 2963 QDFFRBN $T=492280 991320 1 180 $X=480500 $Y=990940
X1503 2967 252 2950 2 1 3026 QDFFRBN $T=480500 1031640 0 0 $X=480500 $Y=1031260
X1504 2977 2637 2970 2 1 2994 QDFFRBN $T=482360 971160 0 0 $X=482360 $Y=970780
X1505 2991 252 309 2 1 2999 QDFFRBN $T=484840 1082040 1 0 $X=484840 $Y=1076620
X1506 3003 253 305 2 1 329 QDFFRBN $T=487940 910680 1 0 $X=487940 $Y=905260
X1507 3009 253 2951 2 1 330 QDFFRBN $T=489180 910680 0 0 $X=489180 $Y=910300
X1508 3036 253 2951 2 1 2974 QDFFRBN $T=500960 930840 0 180 $X=489180 $Y=925420
X1509 3034 2637 2887 2 1 2989 QDFFRBN $T=500960 1021560 1 180 $X=489180 $Y=1021180
X1510 3065 252 2950 2 1 3008 QDFFRBN $T=500960 1041720 1 180 $X=489180 $Y=1041340
X1511 3068 2637 2941 2 1 3013 QDFFRBN $T=504060 951000 1 180 $X=492280 $Y=950620
X1512 3078 2637 2955 2 1 2189 QDFFRBN $T=504060 991320 0 180 $X=492280 $Y=985900
X1513 3066 253 2807 2 1 3021 QDFFRBN $T=505300 940920 0 180 $X=493520 $Y=935500
X1514 3042 2637 2955 2 1 2986 QDFFRBN $T=505300 1001400 1 180 $X=493520 $Y=1001020
X1515 3070 2637 2955 2 1 3020 QDFFRBN $T=505920 991320 1 180 $X=494140 $Y=990940
X1516 3038 253 2951 2 1 317 QDFFRBN $T=506540 920760 0 180 $X=494760 $Y=915340
X1517 3084 2637 2970 2 1 3018 QDFFRBN $T=506540 971160 1 180 $X=494760 $Y=970780
X1518 3032 252 3079 2 1 3083 QDFFRBN $T=494760 1031640 0 0 $X=494760 $Y=1031260
X1519 3092 252 3071 2 1 3002 QDFFRBN $T=508400 1071960 0 180 $X=496620 $Y=1066540
X1520 3081 252 3071 2 1 3057 QDFFRBN $T=509640 1051800 1 180 $X=497860 $Y=1051420
X1521 3119 253 305 2 1 328 QDFFRBN $T=510880 900600 1 180 $X=499100 $Y=900220
X1522 3094 253 2807 2 1 3073 QDFFRBN $T=512120 940920 1 180 $X=500340 $Y=940540
X1523 3058 253 2807 2 1 2584 QDFFRBN $T=502820 930840 1 0 $X=502820 $Y=925420
X1524 3147 252 3071 2 1 337 QDFFRBN $T=516460 1061880 1 180 $X=504680 $Y=1061500
X1525 3148 2637 3115 2 1 3091 QDFFRBN $T=517080 1021560 0 180 $X=505300 $Y=1016140
X1526 3098 252 354 2 1 3125 QDFFRBN $T=505920 1082040 1 0 $X=505920 $Y=1076620
X1527 3102 2637 3144 2 1 358 QDFFRBN $T=506540 991320 0 0 $X=506540 $Y=990940
X1528 3107 253 3134 2 1 3156 QDFFRBN $T=507160 951000 1 0 $X=507160 $Y=945580
X1529 3108 2637 3144 2 1 2509 QDFFRBN $T=507160 971160 0 0 $X=507160 $Y=970780
X1530 3109 2637 3144 2 1 2413 QDFFRBN $T=507160 981240 1 0 $X=507160 $Y=975820
X1531 3111 2637 3134 2 1 2123 QDFFRBN $T=507780 971160 1 0 $X=507780 $Y=965740
X1532 3164 253 2807 2 1 3112 QDFFRBN $T=520180 920760 1 180 $X=508400 $Y=920380
X1533 3170 253 3134 2 1 3099 QDFFRBN $T=520800 930840 1 180 $X=509020 $Y=930460
X1534 3124 2637 3157 2 1 3143 QDFFRBN $T=509640 1011480 1 0 $X=509640 $Y=1006060
X1535 3131 2637 3157 2 1 3117 QDFFRBN $T=510880 1011480 0 0 $X=510880 $Y=1011100
X1536 3133 252 3115 2 1 3189 QDFFRBN $T=511500 1031640 0 0 $X=511500 $Y=1031260
X1537 3138 2637 3134 2 1 2272 QDFFRBN $T=512740 961080 0 0 $X=512740 $Y=960700
X1538 3168 253 357 2 1 349 QDFFRBN $T=526380 900600 1 180 $X=514600 $Y=900220
X1539 3210 2637 3144 2 1 3151 QDFFRBN $T=528240 1001400 1 180 $X=516460 $Y=1001020
X1540 3165 2637 3134 2 1 3188 QDFFRBN $T=518320 961080 1 0 $X=518320 $Y=955660
X1541 3167 252 360 2 1 3207 QDFFRBN $T=518320 1061880 0 0 $X=518320 $Y=1061500
X1542 3172 2637 3144 2 1 366 QDFFRBN $T=520180 991320 0 0 $X=520180 $Y=990940
X1543 3191 2637 3115 2 1 3126 QDFFRBN $T=532580 1021560 1 180 $X=520800 $Y=1021180
X1544 3181 2637 3223 2 1 3199 QDFFRBN $T=521420 981240 1 0 $X=521420 $Y=975820
X1545 3186 253 3228 2 1 3212 QDFFRBN $T=522040 910680 0 0 $X=522040 $Y=910300
X1546 3184 253 3228 2 1 2261 QDFFRBN $T=523280 930840 0 0 $X=523280 $Y=930460
X1547 3204 253 3228 2 1 3178 QDFFRBN $T=523900 920760 0 0 $X=523900 $Y=920380
X1548 3202 2637 3157 2 1 378 QDFFRBN $T=523900 1021560 1 0 $X=523900 $Y=1016140
X1549 3206 252 360 2 1 381 QDFFRBN $T=524520 1071960 1 0 $X=524520 $Y=1066540
X1550 3246 2637 3071 2 1 3174 QDFFRBN $T=537540 1051800 0 180 $X=525760 $Y=1046380
X1551 3267 3257 3223 2 1 3214 QDFFRBN $T=538780 961080 1 180 $X=527000 $Y=960700
X1552 3248 2637 3115 2 1 3171 QDFFRBN $T=539400 1031640 1 180 $X=527620 $Y=1031260
X1553 3273 380 357 2 1 370 QDFFRBN $T=541880 900600 1 180 $X=530100 $Y=900220
X1554 3230 2637 3232 2 1 3284 QDFFRBN $T=530100 1001400 0 0 $X=530100 $Y=1001020
X1555 3251 380 3294 2 1 3330 QDFFRBN $T=534440 940920 1 0 $X=534440 $Y=935500
X1556 3252 2637 3157 2 1 390 QDFFRBN $T=534440 1021560 0 0 $X=534440 $Y=1021180
X1557 3264 3257 3144 2 1 3236 QDFFRBN $T=546840 991320 1 180 $X=535060 $Y=990940
X1558 3256 380 3294 2 1 3318 QDFFRBN $T=535680 910680 0 0 $X=535680 $Y=910300
X1559 3317 3257 3232 2 1 2219 QDFFRBN $T=547460 1031640 0 180 $X=535680 $Y=1026220
X1560 3261 3257 3223 2 1 3315 QDFFRBN $T=536300 981240 1 0 $X=536300 $Y=975820
X1561 3320 399 360 2 1 3260 QDFFRBN $T=548080 1071960 0 180 $X=536300 $Y=1066540
X1562 3278 380 3294 2 1 3275 QDFFRBN $T=538780 920760 0 0 $X=538780 $Y=920380
X1563 3279 3257 3223 2 1 2305 QDFFRBN $T=539400 981240 0 0 $X=539400 $Y=980860
X1564 3281 3257 3307 2 1 3339 QDFFRBN $T=540020 961080 1 0 $X=540020 $Y=955660
X1565 3286 3257 3307 2 1 409 QDFFRBN $T=541260 961080 0 0 $X=541260 $Y=960700
X1566 3302 3257 3232 2 1 2231 QDFFRBN $T=543120 1011480 1 0 $X=543120 $Y=1006060
X1567 3366 3257 3232 2 1 3308 QDFFRBN $T=556140 1001400 1 180 $X=544360 $Y=1001020
X1568 3312 399 3356 2 1 3371 QDFFRBN $T=544360 1061880 1 0 $X=544360 $Y=1056460
X1569 3313 399 360 2 1 3322 QDFFRBN $T=544360 1071960 0 0 $X=544360 $Y=1071580
X1570 3389 380 3258 2 1 3329 QDFFRBN $T=559860 940920 0 180 $X=548080 $Y=935500
X1571 3335 380 3294 2 1 3370 QDFFRBN $T=548700 930840 1 0 $X=548700 $Y=925420
X1572 3380 380 3294 2 1 3285 QDFFRBN $T=561720 910680 1 180 $X=549940 $Y=910300
X1573 3342 3257 3385 2 1 3344 QDFFRBN $T=549940 1031640 1 0 $X=549940 $Y=1026220
X1574 3340 3257 3306 2 1 408 QDFFRBN $T=549940 1041720 1 0 $X=549940 $Y=1036300
X1575 3404 3257 3307 2 1 3355 QDFFRBN $T=564200 971160 1 180 $X=552420 $Y=970780
X1576 3350 3257 3232 2 1 2236 QDFFRBN $T=552420 1021560 0 0 $X=552420 $Y=1021180
X1577 3428 3257 3307 2 1 2674 QDFFRBN $T=567300 961080 1 180 $X=555520 $Y=960700
X1578 3376 3257 3232 2 1 3423 QDFFRBN $T=556140 1021560 1 0 $X=556140 $Y=1016140
X1579 3379 3257 3306 2 1 436 QDFFRBN $T=556760 1041720 0 0 $X=556760 $Y=1041340
X1580 3442 380 3407 2 1 3390 QDFFRBN $T=570400 951000 1 180 $X=558620 $Y=950620
X1581 3394 3257 3385 2 1 3434 QDFFRBN $T=558620 1001400 0 0 $X=558620 $Y=1001020
X1582 3457 380 3397 2 1 2598 QDFFRBN $T=572880 930840 1 180 $X=561100 $Y=930460
X1583 3431 380 3258 2 1 3365 QDFFRBN $T=572880 940920 0 180 $X=561100 $Y=935500
X1584 3444 399 3356 2 1 425 QDFFRBN $T=572880 1061880 1 180 $X=561100 $Y=1061500
X1585 3421 380 3397 2 1 3466 QDFFRBN $T=562960 930840 1 0 $X=562960 $Y=925420
X1586 428 380 3461 2 1 443 QDFFRBN $T=563580 900600 0 0 $X=563580 $Y=900220
X1587 3419 380 3461 2 1 444 QDFFRBN $T=563580 910680 1 0 $X=563580 $Y=905260
X1588 3427 380 3461 2 1 3435 QDFFRBN $T=564200 910680 0 0 $X=564200 $Y=910300
X1589 3439 3257 3385 2 1 429 QDFFRBN $T=575980 1031640 0 180 $X=564200 $Y=1026220
X1590 3433 3257 3473 2 1 3468 QDFFRBN $T=565440 991320 0 0 $X=565440 $Y=990940
X1591 3491 399 3391 2 1 3416 QDFFRBN $T=579080 1051800 0 180 $X=567300 $Y=1046380
X1592 3446 399 447 2 1 3448 QDFFRBN $T=567920 1082040 0 0 $X=567920 $Y=1081660
X1593 3452 3257 3473 2 1 3408 QDFFRBN $T=568540 981240 0 0 $X=568540 $Y=980860
X1594 3450 3257 3306 2 1 440 QDFFRBN $T=568540 1031640 0 0 $X=568540 $Y=1031260
X1595 3488 399 3356 2 1 3412 QDFFRBN $T=580320 1061880 0 180 $X=568540 $Y=1056460
X1596 3453 3257 3385 2 1 445 QDFFRBN $T=569160 1011480 0 0 $X=569160 $Y=1011100
X1597 3447 3257 3407 2 1 3481 QDFFRBN $T=569780 961080 0 0 $X=569780 $Y=960700
X1598 3502 399 3391 2 1 438 QDFFRBN $T=581560 1041720 1 180 $X=569780 $Y=1041340
X1599 3469 3257 3473 2 1 446 QDFFRBN $T=572880 1001400 0 0 $X=572880 $Y=1001020
X1600 3475 399 459 2 1 450 QDFFRBN $T=572880 1071960 0 0 $X=572880 $Y=1071580
X1601 3522 380 3397 2 1 3478 QDFFRBN $T=585900 940920 0 180 $X=574120 $Y=935500
X1602 3479 380 3511 2 1 3529 QDFFRBN $T=574740 930840 0 0 $X=574740 $Y=930460
X1603 3489 380 3397 2 1 3462 QDFFRBN $T=576600 920760 0 0 $X=576600 $Y=920380
X1604 3493 380 3461 2 1 3521 QDFFRBN $T=577840 910680 1 0 $X=577840 $Y=905260
X1605 3545 3257 3473 2 1 3490 QDFFRBN $T=591480 991320 1 180 $X=579700 $Y=990940
X1606 3551 399 3391 2 1 3507 QDFFRBN $T=593340 1051800 0 180 $X=581560 $Y=1046380
X1607 3566 3257 3539 2 1 3510 QDFFRBN $T=595200 1011480 1 180 $X=583420 $Y=1011100
X1608 3530 3257 3559 2 1 3499 QDFFRBN $T=584660 1031640 1 0 $X=584660 $Y=1026220
X1609 3578 380 3407 2 1 471 QDFFRBN $T=597060 951000 0 180 $X=585280 $Y=945580
X1610 3554 399 459 2 1 3527 QDFFRBN $T=597680 1071960 0 180 $X=585900 $Y=1066540
X1611 3542 3257 3539 2 1 3552 QDFFRBN $T=587140 1001400 0 0 $X=587140 $Y=1001020
X1612 3576 380 3511 2 1 3218 QDFFRBN $T=599540 940920 0 180 $X=587760 $Y=935500
X1613 3523 3257 3539 2 1 452 QDFFRBN $T=599540 971160 1 180 $X=587760 $Y=970780
X1614 486 399 459 2 1 474 QDFFRBN $T=600160 1082040 1 180 $X=588380 $Y=1081660
X1615 3574 380 3407 2 1 3546 QDFFRBN $T=600780 961080 0 180 $X=589000 $Y=955660
X1616 3572 3257 3539 2 1 3544 QDFFRBN $T=600780 991320 0 180 $X=589000 $Y=985900
X1617 3605 380 3407 2 1 476 QDFFRBN $T=602020 951000 1 180 $X=590240 $Y=950620
X1618 3549 3257 3582 2 1 3534 QDFFRBN $T=590240 1021560 1 0 $X=590240 $Y=1016140
X1619 3547 399 3356 2 1 467 QDFFRBN $T=602640 1061880 1 180 $X=590860 $Y=1061500
X1620 495 380 3461 2 1 479 QDFFRBN $T=603260 910680 0 180 $X=591480 $Y=905260
X1621 3557 399 3592 2 1 3571 QDFFRBN $T=592100 1051800 0 0 $X=592100 $Y=1051420
X1622 3560 399 459 2 1 3625 QDFFRBN $T=592720 1082040 1 0 $X=592720 $Y=1076620
X1623 3567 3257 3559 2 1 3619 QDFFRBN $T=593960 1041720 1 0 $X=593960 $Y=1036300
X1624 3575 3257 3592 2 1 3641 QDFFRBN $T=595820 1041720 0 0 $X=595820 $Y=1041340
X1625 3579 3257 3539 2 1 505 QDFFRBN $T=597060 981240 1 0 $X=597060 $Y=975820
X1626 3613 380 3511 2 1 2631 QDFFRBN $T=609460 930840 0 180 $X=597680 $Y=925420
X1627 3581 3257 3610 2 1 3650 QDFFRBN $T=597680 991320 0 0 $X=597680 $Y=990940
X1628 3585 3257 3559 2 1 508 QDFFRBN $T=598300 1031640 1 0 $X=598300 $Y=1026220
X1629 3593 3257 3559 2 1 3660 QDFFRBN $T=599540 1031640 0 0 $X=599540 $Y=1031260
X1630 3597 3257 3582 2 1 510 QDFFRBN $T=600160 1001400 1 0 $X=600160 $Y=995980
X1631 3598 3257 3610 2 1 511 QDFFRBN $T=600160 1011480 1 0 $X=600160 $Y=1006060
X1632 3601 380 3511 2 1 478 QDFFRBN $T=600780 930840 0 0 $X=600780 $Y=930460
X1633 3622 3257 3539 2 1 2496 QDFFRBN $T=612560 971160 1 180 $X=600780 $Y=970780
X1634 3632 3257 3610 2 1 481 QDFFRBN $T=613800 991320 0 180 $X=602020 $Y=985900
X1635 3604 3257 3582 2 1 3588 QDFFRBN $T=602020 1021560 1 0 $X=602020 $Y=1016140
X1636 3653 399 3592 2 1 3602 QDFFRBN $T=615040 1071960 0 180 $X=603260 $Y=1066540
X1637 3662 380 499 2 1 3603 QDFFRBN $T=615660 920760 0 180 $X=603880 $Y=915340
X1638 3658 399 3592 2 1 3612 QDFFRBN $T=615660 1061880 1 180 $X=603880 $Y=1061500
X1639 3615 3257 3610 2 1 521 QDFFRBN $T=604500 1011480 0 0 $X=604500 $Y=1011100
X1640 3626 380 499 2 1 3627 QDFFRBN $T=605740 910680 0 0 $X=605740 $Y=910300
X1641 3617 380 3511 2 1 435 QDFFRBN $T=617520 940920 1 180 $X=605740 $Y=940540
X1642 3631 380 3669 2 1 3691 QDFFRBN $T=606360 951000 1 0 $X=606360 $Y=945580
X1643 3635 380 3669 2 1 525 QDFFRBN $T=607600 951000 0 0 $X=607600 $Y=950620
X1644 3642 380 3669 2 1 3487 QDFFRBN $T=608220 961080 1 0 $X=608220 $Y=955660
X1645 3703 3257 3610 2 1 3638 QDFFRBN $T=620000 981240 1 180 $X=608220 $Y=980860
X1646 3698 380 3511 2 1 3589 QDFFRBN $T=621240 930840 0 180 $X=609460 $Y=925420
X1647 3655 3257 3710 2 1 3692 QDFFRBN $T=611320 981240 1 0 $X=611320 $Y=975820
X1648 3667 380 3723 2 1 3728 QDFFRBN $T=613800 940920 1 0 $X=613800 $Y=935500
X1649 3720 3257 3582 2 1 3670 QDFFRBN $T=626200 1021560 0 180 $X=614420 $Y=1016140
X1650 3732 399 527 2 1 3689 QDFFRBN $T=628680 1071960 1 180 $X=616900 $Y=1071580
X1651 3672 3257 3710 2 1 3694 QDFFRBN $T=618140 991320 0 0 $X=618140 $Y=990940
X1652 3705 3257 3753 2 1 535 QDFFRBN $T=618140 1011480 0 0 $X=618140 $Y=1011100
X1653 3707 399 527 2 1 3744 QDFFRBN $T=618140 1071960 1 0 $X=618140 $Y=1066540
X1654 3668 380 499 2 1 3621 QDFFRBN $T=631160 910680 0 180 $X=619380 $Y=905260
X1655 3714 380 3710 2 1 3724 QDFFRBN $T=620000 961080 1 0 $X=620000 $Y=955660
X1656 3749 3257 3710 2 1 3550 QDFFRBN $T=631780 1001400 0 180 $X=620000 $Y=995980
X1657 536 380 499 2 1 524 QDFFRBN $T=632400 900600 1 180 $X=620620 $Y=900220
X1658 3716 380 3723 2 1 2597 QDFFRBN $T=633020 910680 1 180 $X=621240 $Y=910300
X1659 3717 399 3759 2 1 3738 QDFFRBN $T=621240 1041720 0 0 $X=621240 $Y=1041340
X1660 3772 380 3723 2 1 487 QDFFRBN $T=633640 920760 1 180 $X=621860 $Y=920380
X1661 3727 3257 3710 2 1 3569 QDFFRBN $T=621860 981240 0 0 $X=621860 $Y=980860
X1662 3792 380 3723 2 1 531 QDFFRBN $T=635500 930840 0 180 $X=623720 $Y=925420
X1663 3763 3257 3730 2 1 3611 QDFFRBN $T=636120 1021560 1 180 $X=624340 $Y=1021180
X1664 3793 399 3759 2 1 3743 QDFFRBN $T=636120 1051800 0 180 $X=624340 $Y=1046380
X1665 3755 380 3723 2 1 3785 QDFFRBN $T=627440 940920 1 0 $X=627440 $Y=935500
X1666 3775 399 527 2 1 3820 QDFFRBN $T=629920 1082040 1 0 $X=629920 $Y=1076620
X1667 3811 380 3723 2 1 3776 QDFFRBN $T=642320 920760 0 180 $X=630540 $Y=915340
X1668 3779 399 554 2 1 3771 QDFFRBN $T=630540 1071960 1 0 $X=630540 $Y=1066540
X1669 3818 3257 3753 2 1 3766 QDFFRBN $T=642940 1011480 1 180 $X=631160 $Y=1011100
X1670 540 399 554 2 1 547 QDFFRBN $T=631160 1082040 0 0 $X=631160 $Y=1081660
X1671 3787 380 3669 2 1 539 QDFFRBN $T=631780 961080 1 0 $X=631780 $Y=955660
X1672 3784 3257 3794 2 1 550 QDFFRBN $T=631780 1001400 1 0 $X=631780 $Y=995980
X1673 3805 3257 3730 2 1 537 QDFFRBN $T=643560 1021560 0 180 $X=631780 $Y=1016140
X1674 3844 3257 3753 2 1 3790 QDFFRBN $T=645420 1001400 1 180 $X=633640 $Y=1001020
X1675 3804 3257 3730 2 1 3764 QDFFRBN $T=645420 1031640 1 180 $X=633640 $Y=1031260
X1676 3807 399 527 2 1 3791 QDFFRBN $T=645420 1061880 1 180 $X=633640 $Y=1061500
X1677 545 380 3824 2 1 563 QDFFRBN $T=634880 900600 0 0 $X=634880 $Y=900220
X1678 3798 380 3824 2 1 3825 QDFFRBN $T=636120 910680 0 0 $X=636120 $Y=910300
X1679 3800 399 3759 2 1 3829 QDFFRBN $T=636120 1041720 0 0 $X=636120 $Y=1041340
X1680 3809 380 3821 2 1 3865 QDFFRBN $T=638600 930840 1 0 $X=638600 $Y=925420
X1681 3850 3819 3794 2 1 555 QDFFRBN $T=651620 971160 0 180 $X=639840 $Y=965740
X1682 3816 3819 3669 2 1 3599 QDFFRBN $T=640460 951000 0 0 $X=640460 $Y=950620
X1683 3817 3819 3669 2 1 3873 QDFFRBN $T=640460 961080 0 0 $X=640460 $Y=960700
X1684 556 380 3824 2 1 3848 QDFFRBN $T=641080 910680 1 0 $X=641080 $Y=905260
X1685 3835 3257 3874 2 1 3596 QDFFRBN $T=644180 1021560 0 0 $X=644180 $Y=1021180
X1686 3837 399 554 2 1 3855 QDFFRBN $T=644180 1071960 1 0 $X=644180 $Y=1066540
X1687 3842 3257 3874 2 1 3884 QDFFRBN $T=645420 1011480 0 0 $X=645420 $Y=1011100
X1688 3849 399 3890 2 1 3899 QDFFRBN $T=646660 1061880 0 0 $X=646660 $Y=1061500
X1689 3905 3819 3821 2 1 564 QDFFRBN $T=659680 951000 0 180 $X=647900 $Y=945580
X1690 3853 3257 3874 2 1 3607 QDFFRBN $T=647900 1001400 0 0 $X=647900 $Y=1001020
X1691 3856 3819 3901 2 1 3869 QDFFRBN $T=649140 981240 1 0 $X=649140 $Y=975820
X1692 3862 3257 3759 2 1 3828 QDFFRBN $T=660920 1041720 1 180 $X=649140 $Y=1041340
X1693 3861 3819 3901 2 1 3733 QDFFRBN $T=649760 991320 0 0 $X=649760 $Y=990940
X1694 3909 586 3824 2 1 570 QDFFRBN $T=662780 910680 1 180 $X=651000 $Y=910300
X1695 590 399 554 2 1 571 QDFFRBN $T=662780 1082040 1 180 $X=651000 $Y=1081660
X1696 3935 3819 3874 2 1 3880 QDFFRBN $T=665260 1031640 0 180 $X=653480 $Y=1026220
X1697 3886 3257 3874 2 1 581 QDFFRBN $T=654100 1021560 1 0 $X=654100 $Y=1016140
X1698 3974 3819 3903 2 1 3904 QDFFRBN $T=669600 920760 1 180 $X=657820 $Y=920380
X1699 3939 599 3890 2 1 3906 QDFFRBN $T=669600 1071960 0 180 $X=657820 $Y=1066540
X1700 3936 599 3890 2 1 3908 QDFFRBN $T=672080 1061880 1 180 $X=660300 $Y=1061500
X1701 3960 3819 3903 2 1 3883 QDFFRBN $T=672700 930840 0 180 $X=660920 $Y=925420
X1702 3929 586 593 2 1 3945 QDFFRBN $T=661540 920760 1 0 $X=661540 $Y=915340
X1703 3958 3819 3874 2 1 592 QDFFRBN $T=673320 1001400 1 180 $X=661540 $Y=1001020
X1704 595 586 593 2 1 614 QDFFRBN $T=664020 900600 0 0 $X=664020 $Y=900220
X1705 3924 586 593 2 1 3902 QDFFRBN $T=664020 910680 1 0 $X=664020 $Y=905260
X1706 3950 3819 4003 2 1 3609 QDFFRBN $T=664640 940920 1 0 $X=664640 $Y=935500
X1707 3977 3819 3901 2 1 3922 QDFFRBN $T=676420 981240 0 180 $X=664640 $Y=975820
X1708 3953 599 3890 2 1 618 QDFFRBN $T=665260 1061880 1 0 $X=665260 $Y=1056460
X1709 3957 586 4003 2 1 624 QDFFRBN $T=665880 910680 0 0 $X=665880 $Y=910300
X1710 3981 3819 4024 2 1 3934 QDFFRBN $T=668360 1011480 0 0 $X=668360 $Y=1011100
X1711 3967 3819 3972 2 1 3923 QDFFRBN $T=680140 1051800 0 180 $X=668360 $Y=1046380
X1712 4002 3819 3972 2 1 3919 QDFFRBN $T=680760 1041720 0 180 $X=668980 $Y=1036300
X1713 4006 599 3890 2 1 602 QDFFRBN $T=680760 1071960 1 180 $X=668980 $Y=1071580
X1714 3963 3819 3901 2 1 3639 QDFFRBN $T=681380 1011480 0 180 $X=669600 $Y=1006060
X1715 3986 3819 3972 2 1 3978 QDFFRBN $T=682000 1031640 1 180 $X=670220 $Y=1031260
X1716 4056 3819 3901 2 1 4000 QDFFRBN $T=683240 971160 1 180 $X=671460 $Y=970780
X1717 4022 3819 4060 2 1 640 QDFFRBN $T=675800 1021560 1 0 $X=675800 $Y=1016140
X1718 4026 599 4019 2 1 4092 QDFFRBN $T=676420 1071960 1 0 $X=676420 $Y=1066540
X1719 641 586 4003 2 1 619 QDFFRBN $T=688820 900600 1 180 $X=677040 $Y=900220
X1720 4027 3819 4003 2 1 3954 QDFFRBN $T=677660 930840 0 0 $X=677660 $Y=930460
X1721 4101 3819 4058 2 1 3898 QDFFRBN $T=690680 940920 0 180 $X=678900 $Y=935500
X1722 4042 3819 4064 2 1 4108 QDFFRBN $T=678900 981240 1 0 $X=678900 $Y=975820
X1723 4097 3819 4060 2 1 4040 QDFFRBN $T=690680 1021560 1 180 $X=678900 $Y=1021180
X1724 4105 3819 4064 2 1 4043 QDFFRBN $T=691300 991320 1 180 $X=679520 $Y=990940
X1725 4110 3819 4024 2 1 4051 QDFFRBN $T=691920 1001400 1 180 $X=680140 $Y=1001020
X1726 4119 3819 4058 2 1 3993 QDFFRBN $T=693160 951000 0 180 $X=681380 $Y=945580
X1727 4106 3819 4003 2 1 3982 QDFFRBN $T=693780 910680 1 180 $X=682000 $Y=910300
X1728 4068 3819 4064 2 1 4063 QDFFRBN $T=683240 971160 0 0 $X=683240 $Y=970780
X1729 4169 3819 4003 2 1 4048 QDFFRBN $T=699360 930840 0 180 $X=687580 $Y=925420
X1730 4152 3819 4058 2 1 628 QDFFRBN $T=699360 961080 1 180 $X=687580 $Y=960700
X1731 4143 3819 4058 2 1 4095 QDFFRBN $T=699980 951000 1 180 $X=688200 $Y=950620
X1732 4102 3819 4060 2 1 3949 QDFFRBN $T=688820 1021560 1 0 $X=688820 $Y=1016140
X1733 4129 3819 4124 2 1 4009 QDFFRBN $T=701220 1041720 1 180 $X=689440 $Y=1041340
X1734 4107 599 650 2 1 4125 QDFFRBN $T=689440 1082040 1 0 $X=689440 $Y=1076620
X1735 4109 586 651 2 1 4076 QDFFRBN $T=690060 900600 0 0 $X=690060 $Y=900220
X1736 4156 3819 4058 2 1 3851 QDFFRBN $T=702460 940920 1 180 $X=690680 $Y=940540
X1737 4099 599 4019 2 1 4120 QDFFRBN $T=690680 1071960 1 0 $X=690680 $Y=1066540
X1738 4121 599 4019 2 1 3992 QDFFRBN $T=691300 1061880 1 0 $X=691300 $Y=1056460
X1739 4165 3819 4134 2 1 3808 QDFFRBN $T=703700 1001400 0 180 $X=691920 $Y=995980
X1740 4144 3819 4060 2 1 4085 QDFFRBN $T=704320 1021560 1 180 $X=692540 $Y=1021180
X1741 4157 3819 4134 2 1 4127 QDFFRBN $T=704940 991320 1 180 $X=693160 $Y=990940
X1742 4130 3819 4064 2 1 4197 QDFFRBN $T=693780 981240 1 0 $X=693780 $Y=975820
X1743 4182 586 4153 2 1 4140 QDFFRBN $T=708040 910680 1 180 $X=696260 $Y=910300
X1744 4185 3819 4060 2 1 639 QDFFRBN $T=708040 1011480 1 180 $X=696260 $Y=1011100
X1745 4160 3819 4153 2 1 3907 QDFFRBN $T=698740 930840 0 0 $X=698740 $Y=930460
X1746 4162 3819 4153 2 1 4203 QDFFRBN $T=699360 940920 1 0 $X=699360 $Y=935500
X1747 4163 3819 4124 2 1 4148 QDFFRBN $T=699360 1051800 1 0 $X=699360 $Y=1046380
X1748 4172 3819 4064 2 1 4235 QDFFRBN $T=700600 971160 1 0 $X=700600 $Y=965740
X1749 4173 3819 4217 2 1 4238 QDFFRBN $T=700600 1001400 0 0 $X=700600 $Y=1001020
X1750 4186 599 4221 2 1 4052 QDFFRBN $T=702460 1071960 1 0 $X=702460 $Y=1066540
X1751 4187 586 4232 2 1 4147 QDFFRBN $T=703700 900600 0 0 $X=703700 $Y=900220
X1752 4189 599 4221 2 1 4225 QDFFRBN $T=703700 1061880 1 0 $X=703700 $Y=1056460
X1753 4201 3819 4236 2 1 4178 QDFFRBN $T=705560 1041720 1 0 $X=705560 $Y=1036300
X1754 4207 3819 4248 2 1 4252 QDFFRBN $T=706180 951000 1 0 $X=706180 $Y=945580
X1755 4208 3819 4217 2 1 665 QDFFRBN $T=706800 991320 0 0 $X=706800 $Y=990940
X1756 4210 3819 4236 2 1 4194 QDFFRBN $T=706800 1021560 0 0 $X=706800 $Y=1021180
X1757 4212 3819 4253 2 1 4198 QDFFRBN $T=707420 981240 1 0 $X=707420 $Y=975820
X1758 4213 3819 4253 2 1 670 QDFFRBN $T=707420 1011480 1 0 $X=707420 $Y=1006060
X1759 4293 3819 651 2 1 4233 QDFFRBN $T=723540 910680 1 180 $X=711760 $Y=910300
X1760 4257 3819 4248 2 1 4115 QDFFRBN $T=723540 930840 0 180 $X=711760 $Y=925420
X1761 4258 3819 4153 2 1 4223 QDFFRBN $T=724160 940920 0 180 $X=712380 $Y=935500
X1762 4188 3819 4248 2 1 4211 QDFFRBN $T=712380 971160 1 0 $X=712380 $Y=965740
X1763 4239 599 4124 2 1 681 QDFFRBN $T=712380 1051800 0 0 $X=712380 $Y=1051420
X1764 4244 599 4221 2 1 4285 QDFFRBN $T=713000 1061880 0 0 $X=713000 $Y=1061500
X1765 4303 3819 4253 2 1 4224 QDFFRBN $T=726640 981240 1 180 $X=714860 $Y=980860
X1766 4254 3819 4248 2 1 666 QDFFRBN $T=715480 961080 0 0 $X=715480 $Y=960700
X1767 4317 599 4268 2 1 4214 QDFFRBN $T=727880 1071960 0 180 $X=716100 $Y=1066540
X1768 4294 686 675 2 1 664 QDFFRBN $T=728500 900600 1 180 $X=716720 $Y=900220
X1769 4283 4341 4273 2 1 673 QDFFRBN $T=732840 1021560 0 180 $X=721060 $Y=1016140
X1770 4344 4341 4273 2 1 4277 QDFFRBN $T=732840 1021560 1 180 $X=721060 $Y=1021180
X1771 4373 4341 4248 2 1 4301 QDFFRBN $T=736560 930840 1 180 $X=724780 $Y=930460
X1772 4352 4341 4248 2 1 4270 QDFFRBN $T=736560 940920 0 180 $X=724780 $Y=935500
X1773 4379 4341 4332 2 1 4305 QDFFRBN $T=737180 971160 1 180 $X=725400 $Y=970780
X1774 4383 3819 4232 2 1 4309 QDFFRBN $T=737800 910680 1 180 $X=726020 $Y=910300
X1775 4393 4341 4332 2 1 690 QDFFRBN $T=739660 961080 0 180 $X=727880 $Y=955660
X1776 4395 3819 675 2 1 691 QDFFRBN $T=740280 900600 1 180 $X=728500 $Y=900220
X1777 4372 4341 4332 2 1 4334 QDFFRBN $T=741520 981240 1 180 $X=729740 $Y=980860
X1778 4399 4341 4253 2 1 4046 QDFFRBN $T=741520 1011480 0 180 $X=729740 $Y=1006060
X1779 4410 599 4124 2 1 4337 QDFFRBN $T=741520 1071960 0 180 $X=729740 $Y=1066540
X1780 4319 4341 4401 2 1 4333 QDFFRBN $T=731600 1041720 1 0 $X=731600 $Y=1036300
X1781 4374 4341 4405 2 1 687 QDFFRBN $T=734700 951000 0 0 $X=734700 $Y=950620
X1782 4388 4341 4273 2 1 695 QDFFRBN $T=746480 1011480 1 180 $X=734700 $Y=1011100
X1783 4409 4341 4273 2 1 4356 QDFFRBN $T=746480 1021560 0 180 $X=734700 $Y=1016140
X1784 4406 599 4124 2 1 4376 QDFFRBN $T=747100 1051800 0 180 $X=735320 $Y=1046380
X1785 4440 599 4268 2 1 4377 QDFFRBN $T=747100 1061880 0 180 $X=735320 $Y=1056460
X1786 4385 4341 4408 2 1 4266 QDFFRBN $T=736560 991320 0 0 $X=736560 $Y=990940
X1787 4375 4341 4405 2 1 4287 QDFFRBN $T=749580 940920 0 180 $X=737800 $Y=935500
X1788 4407 4341 4401 2 1 4370 QDFFRBN $T=749580 1031640 0 180 $X=737800 $Y=1026220
X1789 4417 4341 4405 2 1 4345 QDFFRBN $T=750200 930840 0 180 $X=738420 $Y=925420
X1790 4411 4341 4405 2 1 4282 QDFFRBN $T=750200 940920 1 180 $X=738420 $Y=940540
X1791 4430 4341 4332 2 1 4320 QDFFRBN $T=750820 981240 0 180 $X=739040 $Y=975820
X1792 4431 4341 4408 2 1 4343 QDFFRBN $T=751440 1001400 0 180 $X=739660 $Y=995980
X1793 4416 599 4268 2 1 4364 QDFFRBN $T=752680 1082040 0 180 $X=740900 $Y=1076620
X1794 4412 4341 4401 2 1 724 QDFFRBN $T=742140 1021560 0 0 $X=742140 $Y=1021180
X1795 4435 599 4268 2 1 4386 QDFFRBN $T=755160 1071960 0 180 $X=743380 $Y=1066540
X1796 4420 4341 4405 2 1 4335 QDFFRBN $T=755780 910680 1 180 $X=744000 $Y=910300
X1797 4428 599 4401 2 1 697 QDFFRBN $T=755780 1041720 0 180 $X=744000 $Y=1036300
X1798 4474 599 716 2 1 714 QDFFRBN $T=756400 1082040 1 180 $X=744620 $Y=1081660
X1799 4426 4341 4466 2 1 4463 QDFFRBN $T=745860 951000 1 0 $X=745860 $Y=945580
X1800 4427 4341 4459 2 1 4456 QDFFRBN $T=745860 991320 1 0 $X=745860 $Y=985900
X1801 4414 686 4405 2 1 4394 QDFFRBN $T=758260 910680 0 180 $X=746480 $Y=905260
X1802 4429 4341 4466 2 1 4484 QDFFRBN $T=746480 951000 0 0 $X=746480 $Y=950620
X1803 4433 4341 4476 2 1 703 QDFFRBN $T=747720 920760 1 0 $X=747720 $Y=915340
X1804 4436 4341 4478 2 1 4448 QDFFRBN $T=748340 981240 0 0 $X=748340 $Y=980860
X1805 4438 4341 4459 2 1 4487 QDFFRBN $T=748960 1011480 0 0 $X=748960 $Y=1011100
X1806 4439 599 4482 2 1 4501 QDFFRBN $T=748960 1051800 1 0 $X=748960 $Y=1046380
X1807 4443 599 4482 2 1 4502 QDFFRBN $T=749580 1061880 1 0 $X=749580 $Y=1056460
X1808 4451 599 4401 2 1 730 QDFFRBN $T=750820 1031640 0 0 $X=750820 $Y=1031260
X1809 4453 4341 4401 2 1 4516 QDFFRBN $T=751440 1031640 1 0 $X=751440 $Y=1026220
X1810 4457 4341 4459 2 1 4424 QDFFRBN $T=752060 1001400 1 0 $X=752060 $Y=995980
X1811 4468 4341 4476 2 1 4504 QDFFRBN $T=753300 930840 1 0 $X=753300 $Y=925420
X1812 4465 4341 4466 2 1 733 QDFFRBN $T=753300 971160 1 0 $X=753300 $Y=965740
X1813 4467 599 4482 2 1 734 QDFFRBN $T=753300 1051800 0 0 $X=753300 $Y=1051420
X1814 4469 4341 4466 2 1 4525 QDFFRBN $T=753920 961080 0 0 $X=753920 $Y=960700
X1815 4470 4341 4511 2 1 4526 QDFFRBN $T=753920 1021560 0 0 $X=753920 $Y=1021180
X1816 4471 599 731 2 1 4483 QDFFRBN $T=753920 1061880 0 0 $X=753920 $Y=1061500
X1817 4472 4341 4466 2 1 4506 QDFFRBN $T=754540 961080 1 0 $X=754540 $Y=955660
X1818 4475 4341 4476 2 1 4486 QDFFRBN $T=755160 930840 0 0 $X=755160 $Y=930460
X1819 4479 4341 4524 2 1 4460 QDFFRBN $T=756400 910680 0 0 $X=756400 $Y=910300
X1820 4480 4341 4511 2 1 4541 QDFFRBN $T=756400 1021560 1 0 $X=756400 $Y=1016140
X1821 4488 599 740 2 1 4512 QDFFRBN $T=758260 1082040 0 0 $X=758260 $Y=1081660
X1822 4503 4341 4476 2 1 751 QDFFRBN $T=760740 951000 1 0 $X=760740 $Y=945580
X1823 4508 4341 4524 2 1 757 QDFFRBN $T=761360 920760 1 0 $X=761360 $Y=915340
X1824 4499 4341 4478 2 1 4012 QDFFRBN $T=762600 981240 0 0 $X=762600 $Y=980860
X1825 4527 4341 4478 2 1 756 QDFFRBN $T=765080 1001400 1 0 $X=765080 $Y=995980
X1826 4515 4341 4478 2 1 746 QDFFRBN $T=765700 991320 1 0 $X=765700 $Y=985900
X1827 4536 4341 4476 2 1 760 QDFFRBN $T=766940 930840 1 0 $X=766940 $Y=925420
X1828 4537 599 4511 2 1 4585 QDFFRBN $T=766940 1041720 1 0 $X=766940 $Y=1036300
X1829 4552 599 4511 2 1 4510 QDFFRBN $T=769420 1021560 0 0 $X=769420 $Y=1021180
X1830 4563 599 731 2 1 745 QDFFRBN $T=783060 1082040 1 180 $X=771280 $Y=1081660
X1831 4567 4341 4524 2 1 4610 QDFFRBN $T=772520 910680 1 0 $X=772520 $Y=905260
X1832 4589 599 4604 2 1 4580 QDFFRBN $T=784920 1061880 0 180 $X=773140 $Y=1056460
X1833 4595 4341 4524 2 1 4648 QDFFRBN $T=775000 920760 1 0 $X=775000 $Y=915340
X1834 4596 4341 4620 2 1 4654 QDFFRBN $T=775000 951000 1 0 $X=775000 $Y=945580
X1835 4570 599 4604 2 1 744 QDFFRBN $T=786780 1071960 0 180 $X=775000 $Y=1066540
X1836 4669 599 4604 2 1 4605 QDFFRBN $T=788020 1071960 1 180 $X=776240 $Y=1071580
X1837 4626 4341 4620 2 1 4492 QDFFRBN $T=788640 951000 1 180 $X=776860 $Y=950620
X1838 4683 4341 4621 2 1 4617 QDFFRBN $T=790500 981240 0 180 $X=778720 $Y=975820
X1839 4674 4341 4478 2 1 4612 QDFFRBN $T=790500 1001400 0 180 $X=778720 $Y=995980
X1840 4643 4341 4621 2 1 762 QDFFRBN $T=791120 961080 1 180 $X=779340 $Y=960700
X1841 4615 4341 4511 2 1 4622 QDFFRBN $T=791740 1021560 0 180 $X=779960 $Y=1016140
X1842 4629 4341 4621 2 1 4625 QDFFRBN $T=780580 971160 0 0 $X=780580 $Y=970780
X1843 4660 4341 4621 2 1 4581 QDFFRBN $T=793600 991320 0 180 $X=781820 $Y=985900
X1844 4645 4341 4620 2 1 797 QDFFRBN $T=783060 930840 0 0 $X=783060 $Y=930460
X1845 4722 686 784 2 1 778 QDFFRBN $T=797320 900600 1 180 $X=785540 $Y=900220
X1846 4662 4341 4620 2 1 802 QDFFRBN $T=787400 930840 1 0 $X=787400 $Y=925420
X1847 4670 599 804 2 1 793 QDFFRBN $T=787400 1082040 0 0 $X=787400 $Y=1081660
X1848 4691 4341 4692 2 1 4769 QDFFRBN $T=789880 951000 0 0 $X=789880 $Y=950620
X1849 4764 4341 4478 2 1 4689 QDFFRBN $T=801660 1001400 1 180 $X=789880 $Y=1001020
X1850 4642 4341 4708 2 1 4656 QDFFRBN $T=803520 1021560 0 180 $X=791740 $Y=1016140
X1851 4704 4341 4692 2 1 4786 QDFFRBN $T=792360 940920 0 0 $X=792360 $Y=940540
X1852 4707 799 4708 2 1 4696 QDFFRBN $T=792360 1031640 0 0 $X=792360 $Y=1031260
X1853 4712 4341 4621 2 1 4713 QDFFRBN $T=792980 981240 1 0 $X=792980 $Y=975820
X1854 4721 799 4708 2 1 4793 QDFFRBN $T=793600 1031640 1 0 $X=793600 $Y=1026220
X1855 4725 4341 4778 2 1 4514 QDFFRBN $T=794220 1001400 1 0 $X=794220 $Y=995980
X1856 4744 4341 4719 2 1 4554 QDFFRBN $T=797320 930840 0 0 $X=797320 $Y=930460
X1857 4810 686 784 2 1 4760 QDFFRBN $T=811580 900600 1 180 $X=799800 $Y=900220
X1858 4754 4341 4781 2 1 4549 QDFFRBN $T=811580 971160 0 180 $X=799800 $Y=965740
X1859 4767 4341 4719 2 1 813 QDFFRBN $T=812200 920760 1 180 $X=800420 $Y=920380
X1860 4768 799 4708 2 1 4800 QDFFRBN $T=800420 1061880 0 0 $X=800420 $Y=1061500
X1861 4846 4341 4719 2 1 4772 QDFFRBN $T=813440 920760 0 180 $X=801660 $Y=915340
X1862 4776 799 4708 2 1 4822 QDFFRBN $T=801660 1051800 1 0 $X=801660 $Y=1046380
X1863 4759 799 4766 2 1 826 QDFFRBN $T=801660 1071960 1 0 $X=801660 $Y=1066540
X1864 4774 4341 4719 2 1 4847 QDFFRBN $T=802900 930840 1 0 $X=802900 $Y=925420
X1865 4802 799 4856 2 1 4734 QDFFRBN $T=805380 1031640 1 0 $X=805380 $Y=1026220
X1866 4862 4870 4778 2 1 4784 QDFFRBN $T=817780 1001400 0 180 $X=806000 $Y=995980
X1867 4807 4870 4781 2 1 4517 QDFFRBN $T=820260 961080 0 180 $X=808480 $Y=955660
X1868 4857 4870 4909 2 1 4839 QDFFRBN $T=814060 981240 0 0 $X=814060 $Y=980860
X1869 4867 799 4766 2 1 4859 QDFFRBN $T=825840 1061880 1 180 $X=814060 $Y=1061500
X1870 4917 799 4766 2 1 4860 QDFFRBN $T=825840 1071960 1 180 $X=814060 $Y=1071580
X1871 4891 4870 4778 2 1 4863 QDFFRBN $T=826460 1001400 1 180 $X=814680 $Y=1001020
X1872 4921 799 4766 2 1 4873 QDFFRBN $T=827080 1051800 0 180 $X=815300 $Y=1046380
X1873 4913 686 4719 2 1 4874 QDFFRBN $T=827700 920760 1 180 $X=815920 $Y=920380
X1874 4875 686 4914 2 1 4901 QDFFRBN $T=815920 930840 1 0 $X=815920 $Y=925420
X1875 4876 4870 4909 2 1 4818 QDFFRBN $T=815920 981240 1 0 $X=815920 $Y=975820
X1876 4925 686 784 2 1 4879 QDFFRBN $T=828940 900600 1 180 $X=817160 $Y=900220
X1877 4882 4870 4909 2 1 4845 QDFFRBN $T=817160 971160 0 0 $X=817160 $Y=970780
X1878 4940 4870 4908 2 1 4676 QDFFRBN $T=832040 951000 1 180 $X=820260 $Y=950620
X1879 4898 4870 4935 2 1 4946 QDFFRBN $T=820880 991320 1 0 $X=820880 $Y=985900
X1880 4899 799 4856 2 1 4886 QDFFRBN $T=820880 1031640 1 0 $X=820880 $Y=1026220
X1881 4912 4870 4935 2 1 4972 QDFFRBN $T=822740 991320 0 0 $X=822740 $Y=990940
X1882 4979 4870 4908 2 1 4649 QDFFRBN $T=838860 940920 1 180 $X=827080 $Y=940540
X1883 4928 4870 4909 2 1 4974 QDFFRBN $T=827080 971160 1 0 $X=827080 $Y=965740
X1884 4929 799 862 2 1 865 QDFFRBN $T=827080 1082040 0 0 $X=827080 $Y=1081660
X1885 4938 799 4951 2 1 4915 QDFFRBN $T=840100 1071960 1 180 $X=828320 $Y=1071580
X1886 4939 686 4914 2 1 5003 QDFFRBN $T=828940 920760 1 0 $X=828940 $Y=915340
X1887 4920 799 4856 2 1 4904 QDFFRBN $T=840720 1031640 1 180 $X=828940 $Y=1031260
X1888 4943 4870 4908 2 1 4750 QDFFRBN $T=829560 961080 1 0 $X=829560 $Y=955660
X1889 4988 4870 4935 2 1 4941 QDFFRBN $T=841340 981240 0 180 $X=829560 $Y=975820
X1890 4969 799 4856 2 1 852 QDFFRBN $T=841340 1041720 0 180 $X=829560 $Y=1036300
X1891 4996 869 784 2 1 858 QDFFRBN $T=841960 900600 1 180 $X=830180 $Y=900220
X1892 4963 869 4914 2 1 4922 QDFFRBN $T=841960 930840 0 180 $X=830180 $Y=925420
X1893 4958 799 4951 2 1 848 QDFFRBN $T=841960 1071960 0 180 $X=830180 $Y=1066540
X1894 4936 4870 4942 2 1 4947 QDFFRBN $T=830800 1001400 0 0 $X=830800 $Y=1001020
X1895 4948 4870 4942 2 1 4976 QDFFRBN $T=830800 1011480 1 0 $X=830800 $Y=1006060
X1896 4970 799 4951 2 1 4916 QDFFRBN $T=845060 1061880 0 180 $X=833280 $Y=1056460
X1897 4965 799 4856 2 1 4903 QDFFRBN $T=846920 1031640 0 180 $X=835140 $Y=1026220
X1898 4975 799 862 2 1 5036 QDFFRBN $T=835760 1061880 0 0 $X=835760 $Y=1061500
X1899 4985 799 5031 2 1 5005 QDFFRBN $T=837000 1051800 1 0 $X=837000 $Y=1046380
X1900 5002 799 5031 2 1 5068 QDFFRBN $T=840720 1031640 0 0 $X=840720 $Y=1031260
X1901 5008 869 4914 2 1 5048 QDFFRBN $T=841960 920760 0 0 $X=841960 $Y=920380
X1902 5073 4870 4914 2 1 5001 QDFFRBN $T=854360 940920 0 180 $X=842580 $Y=935500
X1903 5011 4870 4935 2 1 5074 QDFFRBN $T=842580 971160 1 0 $X=842580 $Y=965740
X1904 5012 799 5063 2 1 5072 QDFFRBN $T=842580 1021560 0 0 $X=842580 $Y=1021180
X1905 5013 799 5031 2 1 885 QDFFRBN $T=842580 1071960 0 0 $X=842580 $Y=1071580
X1906 5024 869 882 2 1 5078 QDFFRBN $T=843200 910680 1 0 $X=843200 $Y=905260
X1907 5016 4870 5067 2 1 4783 QDFFRBN $T=843200 961080 1 0 $X=843200 $Y=955660
X1908 5025 869 882 2 1 5083 QDFFRBN $T=843820 900600 0 0 $X=843820 $Y=900220
X1909 5022 4870 5063 2 1 5045 QDFFRBN $T=845060 1011480 1 0 $X=845060 $Y=1006060
X1910 5033 4870 5063 2 1 5100 QDFFRBN $T=845680 991320 0 0 $X=845680 $Y=990940
X1911 5038 4870 5067 2 1 5104 QDFFRBN $T=846300 951000 0 0 $X=846300 $Y=950620
X1912 5060 4870 5067 2 1 896 QDFFRBN $T=850020 930840 1 0 $X=850020 $Y=925420
X1913 5061 799 5064 2 1 5069 QDFFRBN $T=850020 1051800 1 0 $X=850020 $Y=1046380
X1914 5134 799 5031 2 1 5088 QDFFRBN $T=866760 1031640 1 180 $X=854980 $Y=1031260
X1915 5151 4870 5067 2 1 5091 QDFFRBN $T=867380 940920 0 180 $X=855600 $Y=935500
X1916 5093 4870 5140 2 1 5137 QDFFRBN $T=856220 961080 1 0 $X=856220 $Y=955660
X1917 5096 799 5143 2 1 5155 QDFFRBN $T=856220 1041720 0 0 $X=856220 $Y=1041340
X1918 5160 869 882 2 1 888 QDFFRBN $T=868620 900600 1 180 $X=856840 $Y=900220
X1919 5103 4870 5140 2 1 5130 QDFFRBN $T=856840 981240 1 0 $X=856840 $Y=975820
X1920 5105 4870 5132 2 1 5128 QDFFRBN $T=858080 981240 0 0 $X=858080 $Y=980860
X1921 5111 4870 5063 2 1 5094 QDFFRBN $T=858700 1011480 1 0 $X=858700 $Y=1006060
X1922 5117 4870 5063 2 1 5185 QDFFRBN $T=859940 1001400 0 0 $X=859940 $Y=1001020
X1923 5189 799 5143 2 1 5123 QDFFRBN $T=873580 1051800 1 180 $X=861800 $Y=1051420
X1924 5164 869 882 2 1 891 QDFFRBN $T=874200 910680 1 180 $X=862420 $Y=910300
X1925 5145 869 5067 2 1 4960 QDFFRBN $T=874200 930840 0 180 $X=862420 $Y=925420
X1926 5139 799 905 2 1 5154 QDFFRBN $T=863660 1071960 0 0 $X=863660 $Y=1071580
X1927 5207 799 905 2 1 5136 QDFFRBN $T=876060 1082040 1 180 $X=864280 $Y=1081660
X1928 5153 869 5200 2 1 5209 QDFFRBN $T=866140 920760 0 0 $X=866140 $Y=920380
X1929 5157 4870 5132 2 1 5202 QDFFRBN $T=866140 991320 1 0 $X=866140 $Y=985900
X1930 5163 4870 5200 2 1 5175 QDFFRBN $T=867380 940920 0 0 $X=867380 $Y=940540
X1931 5152 4870 5140 2 1 914 QDFFRBN $T=868000 971160 0 0 $X=868000 $Y=970780
X1932 5195 4870 5132 2 1 4953 QDFFRBN $T=879780 1011480 1 180 $X=868000 $Y=1011100
X1933 5167 799 5204 2 1 5192 QDFFRBN $T=868000 1031640 1 0 $X=868000 $Y=1026220
X1934 5165 4870 5140 2 1 5221 QDFFRBN $T=869240 961080 1 0 $X=869240 $Y=955660
X1935 907 869 882 2 1 919 QDFFRBN $T=869860 900600 0 0 $X=869860 $Y=900220
X1936 5186 799 5143 2 1 5235 QDFFRBN $T=871100 1041720 0 0 $X=871100 $Y=1041340
X1937 5252 4870 5132 2 1 5187 QDFFRBN $T=883500 1011480 0 180 $X=871720 $Y=1006060
X1938 5188 799 5143 2 1 5199 QDFFRBN $T=871720 1051800 1 0 $X=871720 $Y=1046380
X1939 5241 4870 5200 2 1 5193 QDFFRBN $T=885360 940920 0 180 $X=873580 $Y=935500
X1940 5247 4870 5196 2 1 5171 QDFFRBN $T=885360 981240 0 180 $X=873580 $Y=975820
X1941 5272 4870 5132 2 1 5203 QDFFRBN $T=885980 1001400 0 180 $X=874200 $Y=995980
X1942 5216 799 5265 2 1 5244 QDFFRBN $T=875440 1061880 1 0 $X=875440 $Y=1056460
X1943 5218 799 905 2 1 5253 QDFFRBN $T=876060 1071960 0 0 $X=876060 $Y=1071580
X1944 5261 4870 5200 2 1 5222 QDFFRBN $T=888460 930840 0 180 $X=876680 $Y=925420
X1945 5246 4870 5287 2 1 5281 QDFFRBN $T=881020 951000 1 0 $X=881020 $Y=945580
X1946 5312 4870 5204 2 1 5243 QDFFRBN $T=892800 1031640 0 180 $X=881020 $Y=1026220
X1947 5256 4870 5287 2 1 5330 QDFFRBN $T=882260 961080 0 0 $X=882260 $Y=960700
X1948 5332 5328 5287 2 1 5268 QDFFRBN $T=895900 981240 1 180 $X=884120 $Y=980860
X1949 5282 4870 5287 2 1 5290 QDFFRBN $T=885360 971160 1 0 $X=885360 $Y=965740
X1950 5316 5328 5143 2 1 922 QDFFRBN $T=897760 1041720 1 180 $X=885980 $Y=1041340
X1951 5293 4870 5340 2 1 939 QDFFRBN $T=887220 981240 1 0 $X=887220 $Y=975820
X1952 5286 4870 5321 2 1 942 QDFFRBN $T=888460 930840 0 0 $X=888460 $Y=930460
X1953 5361 4870 5321 2 1 932 QDFFRBN $T=900240 940920 0 180 $X=888460 $Y=935500
X1954 5344 869 937 2 1 5302 QDFFRBN $T=901480 910680 0 180 $X=889700 $Y=905260
X1955 5308 4870 5321 2 1 5311 QDFFRBN $T=889700 920760 0 0 $X=889700 $Y=920380
X1956 5310 799 5265 2 1 5351 QDFFRBN $T=889700 1061880 1 0 $X=889700 $Y=1056460
X1957 5366 946 938 2 1 927 QDFFRBN $T=901480 1071960 1 180 $X=889700 $Y=1071580
X1958 5362 4870 5321 2 1 5299 QDFFRBN $T=902720 930840 0 180 $X=890940 $Y=925420
X1959 5288 5328 5265 2 1 5320 QDFFRBN $T=903960 1031640 1 180 $X=892180 $Y=1031260
X1960 5319 946 938 2 1 5276 QDFFRBN $T=903960 1082040 0 180 $X=892180 $Y=1076620
X1961 5336 4870 5265 2 1 5325 QDFFRBN $T=894040 1031640 1 0 $X=894040 $Y=1026220
X1962 5335 946 938 2 1 5298 QDFFRBN $T=907680 1071960 0 180 $X=895900 $Y=1066540
X1963 5355 4870 5391 2 1 5397 QDFFRBN $T=897760 961080 0 0 $X=897760 $Y=960700
X1964 5346 5328 5333 2 1 5327 QDFFRBN $T=910160 1011480 0 180 $X=898380 $Y=1006060
X1965 5358 5328 5333 2 1 940 QDFFRBN $T=910780 1001400 0 180 $X=899000 $Y=995980
X1966 5365 5328 5340 2 1 5377 QDFFRBN $T=899620 991320 1 0 $X=899620 $Y=985900
X1967 5368 4870 5391 2 1 957 QDFFRBN $T=900240 951000 1 0 $X=900240 $Y=945580
X1968 5364 5328 5340 2 1 5413 QDFFRBN $T=900240 981240 0 0 $X=900240 $Y=980860
X1969 5387 5328 5265 2 1 5309 QDFFRBN $T=912640 1041720 1 180 $X=900860 $Y=1041340
X1970 5381 946 5406 2 1 5427 QDFFRBN $T=902720 1051800 0 0 $X=902720 $Y=1051420
X1971 5382 946 5406 2 1 5424 QDFFRBN $T=902720 1061880 0 0 $X=902720 $Y=1061500
X1972 5373 869 5321 2 1 5370 QDFFRBN $T=915740 920760 1 180 $X=903960 $Y=920380
X1973 5385 5328 5333 2 1 5367 QDFFRBN $T=916980 1011480 1 180 $X=905200 $Y=1011100
X1974 5386 5328 5333 2 1 950 QDFFRBN $T=917600 1021560 0 180 $X=905820 $Y=1016140
X1975 5421 5328 5333 2 1 951 QDFFRBN $T=917600 1021560 1 180 $X=905820 $Y=1021180
X1976 5398 5328 5265 2 1 5443 QDFFRBN $T=906440 1051800 1 0 $X=906440 $Y=1046380
X1977 5430 869 5399 2 1 5345 QDFFRBN $T=918840 940920 0 180 $X=907060 $Y=935500
X1978 5404 5328 5432 2 1 977 QDFFRBN $T=907060 1041720 1 0 $X=907060 $Y=1036300
X1979 5438 973 5391 2 1 5383 QDFFRBN $T=920080 951000 1 180 $X=908300 $Y=950620
X1980 5405 869 974 2 1 5305 QDFFRBN $T=909540 910680 0 0 $X=909540 $Y=910300
X1981 5431 973 5391 2 1 5375 QDFFRBN $T=921320 961080 1 180 $X=909540 $Y=960700
X1982 5409 869 5399 2 1 5472 QDFFRBN $T=910160 930840 1 0 $X=910160 $Y=925420
X1983 5411 946 5406 2 1 994 QDFFRBN $T=910160 1071960 1 0 $X=910160 $Y=1066540
X1984 5414 869 974 2 1 960 QDFFRBN $T=910780 900600 0 0 $X=910780 $Y=900220
X1985 5418 869 5446 2 1 5380 QDFFRBN $T=911400 920760 1 0 $X=911400 $Y=915340
X1986 5455 946 5406 2 1 5412 QDFFRBN $T=923180 1071960 1 180 $X=911400 $Y=1071580
X1987 5439 5328 5432 2 1 966 QDFFRBN $T=923800 1001400 1 180 $X=912020 $Y=1001020
X1988 5419 5328 5451 2 1 986 QDFFRBN $T=912020 1011480 1 0 $X=912020 $Y=1006060
X1989 5469 5328 5204 2 1 965 QDFFRBN $T=923800 1031640 0 180 $X=912020 $Y=1026220
X1990 5437 5328 5432 2 1 5417 QDFFRBN $T=926280 991320 0 180 $X=914500 $Y=985900
X1991 5462 5328 5340 2 1 5393 QDFFRBN $T=927520 981240 0 180 $X=915740 $Y=975820
X1992 5436 973 5487 2 1 5450 QDFFRBN $T=916360 971160 1 0 $X=916360 $Y=965740
X1993 5440 5328 5451 2 1 5504 QDFFRBN $T=917600 1011480 0 0 $X=917600 $Y=1011100
X1994 5449 5328 5451 2 1 5522 QDFFRBN $T=919460 1021560 1 0 $X=919460 $Y=1016140
X1995 5473 869 5446 2 1 5512 QDFFRBN $T=922560 930840 0 0 $X=922560 $Y=930460
X1996 5464 5328 5487 2 1 5423 QDFFRBN $T=934340 981240 1 180 $X=922560 $Y=980860
X1997 5478 973 974 2 1 5544 QDFFRBN $T=923180 910680 1 0 $X=923180 $Y=905260
X1998 5479 973 974 2 1 1010 QDFFRBN $T=923180 910680 0 0 $X=923180 $Y=910300
X1999 5524 973 5446 2 1 5484 QDFFRBN $T=936200 920760 0 180 $X=924420 $Y=915340
X2000 5493 946 5532 2 1 5515 QDFFRBN $T=925040 1051800 0 0 $X=925040 $Y=1051420
X2001 5509 946 5406 2 1 5483 QDFFRBN $T=936820 1071960 1 180 $X=925040 $Y=1071580
X2002 5549 5328 5503 2 1 990 QDFFRBN $T=937440 1001400 1 180 $X=925660 $Y=1001020
X2003 5489 5328 5532 2 1 5447 QDFFRBN $T=925660 1041720 1 0 $X=925660 $Y=1036300
X2004 5502 5328 5503 2 1 5539 QDFFRBN $T=927520 991320 0 0 $X=927520 $Y=990940
X2005 5564 946 5406 2 1 5501 QDFFRBN $T=939300 1071960 0 180 $X=927520 $Y=1066540
X2006 5510 5328 5487 2 1 5520 QDFFRBN $T=929380 971160 1 0 $X=929380 $Y=965740
X2007 5517 5328 5487 2 1 1014 QDFFRBN $T=930620 981240 1 0 $X=930620 $Y=975820
X2008 5547 973 1023 2 1 5612 QDFFRBN $T=935580 910680 0 0 $X=935580 $Y=910300
X2009 5551 5328 5532 2 1 5488 QDFFRBN $T=936200 1031640 1 0 $X=936200 $Y=1026220
X2010 5557 5328 5560 2 1 5641 QDFFRBN $T=936820 1051800 1 0 $X=936820 $Y=1046380
X2011 5563 5328 5503 2 1 5602 QDFFRBN $T=937440 1001400 0 0 $X=937440 $Y=1001020
X2012 5570 5328 5532 2 1 5561 QDFFRBN $T=938680 1021560 0 0 $X=938680 $Y=1021180
X2013 5617 946 1022 2 1 1015 QDFFRBN $T=950460 1071960 1 180 $X=938680 $Y=1071580
X2014 5581 973 5446 2 1 5491 QDFFRBN $T=951080 920760 1 180 $X=939300 $Y=920380
X2015 5578 5328 5503 2 1 5629 QDFFRBN $T=939300 991320 0 0 $X=939300 $Y=990940
X2016 5579 5328 5560 2 1 1032 QDFFRBN $T=939920 1041720 1 0 $X=939920 $Y=1036300
X2017 5583 946 1022 2 1 5623 QDFFRBN $T=940540 1071960 1 0 $X=940540 $Y=1066540
X2018 5619 973 5589 2 1 5582 QDFFRBN $T=953560 971160 0 180 $X=941780 $Y=965740
X2019 5634 973 5446 2 1 5590 QDFFRBN $T=954180 930840 0 180 $X=942400 $Y=925420
X2020 5593 973 5589 2 1 5569 QDFFRBN $T=942400 940920 0 0 $X=942400 $Y=940540
X2021 5599 946 5560 2 1 1008 QDFFRBN $T=954180 1051800 1 180 $X=942400 $Y=1051420
X2022 5600 5328 5589 2 1 5592 QDFFRBN $T=956660 981240 0 180 $X=944880 $Y=975820
X2023 5624 973 5652 2 1 5616 QDFFRBN $T=947360 910680 1 0 $X=947360 $Y=905260
X2024 5628 5328 5503 2 1 5507 QDFFRBN $T=947980 981240 0 0 $X=947980 $Y=980860
X2025 5630 946 1022 2 1 5677 QDFFRBN $T=947980 1082040 0 0 $X=947980 $Y=1081660
X2026 5689 973 5652 2 1 5631 QDFFRBN $T=960380 920760 0 180 $X=948600 $Y=915340
X2027 5679 5328 5503 2 1 5638 QDFFRBN $T=961000 1001400 1 180 $X=949220 $Y=1001020
X2028 5680 946 5560 2 1 5639 QDFFRBN $T=961000 1041720 1 180 $X=949220 $Y=1041340
X2029 5648 5328 5532 2 1 5626 QDFFRBN $T=962240 1021560 1 180 $X=950460 $Y=1021180
X2030 5715 5328 5532 2 1 5658 QDFFRBN $T=964100 1021560 0 180 $X=952320 $Y=1016140
X2031 5645 973 5589 2 1 5672 QDFFRBN $T=952940 951000 1 0 $X=952940 $Y=945580
X2032 5700 973 5682 2 1 5660 QDFFRBN $T=965960 930840 0 180 $X=954180 $Y=925420
X2033 5666 973 5589 2 1 5615 QDFFRBN $T=954800 971160 1 0 $X=954800 $Y=965740
X2034 5675 946 5560 2 1 1027 QDFFRBN $T=956040 1051800 0 0 $X=956040 $Y=1051420
X2035 5737 5328 5697 2 1 5556 QDFFRBN $T=968440 1001400 0 180 $X=956660 $Y=995980
X2036 5686 973 5732 2 1 5724 QDFFRBN $T=957900 961080 0 0 $X=957900 $Y=960700
X2037 5694 5328 5732 2 1 1046 QDFFRBN $T=959140 981240 1 0 $X=959140 $Y=975820
X2038 5703 973 5652 2 1 5681 QDFFRBN $T=960380 910680 0 0 $X=960380 $Y=910300
X2039 5705 973 5652 2 1 5710 QDFFRBN $T=960380 920760 1 0 $X=960380 $Y=915340
X2040 5754 5328 5719 2 1 5684 QDFFRBN $T=972780 1001400 1 180 $X=961000 $Y=1001020
X2041 5673 5328 5697 2 1 5685 QDFFRBN $T=973400 981240 1 180 $X=961620 $Y=980860
X2042 5772 946 5743 2 1 5722 QDFFRBN $T=976500 1041720 1 180 $X=964720 $Y=1041340
X2043 5773 946 1065 2 1 5699 QDFFRBN $T=978980 1082040 0 180 $X=967200 $Y=1076620
X2044 5747 946 1065 2 1 5730 QDFFRBN $T=980220 1071960 1 180 $X=968440 $Y=1071580
X2045 5753 946 5743 2 1 1053 QDFFRBN $T=981460 1051800 1 180 $X=969680 $Y=1051420
X2046 5798 946 5763 2 1 5725 QDFFRBN $T=982080 1061880 0 180 $X=970300 $Y=1056460
X2047 5760 973 5732 2 1 5786 QDFFRBN $T=971540 961080 1 0 $X=971540 $Y=955660
X2048 5792 973 5765 2 1 5741 QDFFRBN $T=985180 920760 0 180 $X=973400 $Y=915340
X2049 5770 973 5682 2 1 1068 QDFFRBN $T=985180 920760 1 180 $X=973400 $Y=920380
X2050 5794 973 5732 2 1 5767 QDFFRBN $T=985800 971160 0 180 $X=974020 $Y=965740
X2051 5811 5328 5732 2 1 5768 QDFFRBN $T=985800 981240 1 180 $X=974020 $Y=980860
X2052 5807 5328 5697 2 1 5647 QDFFRBN $T=985800 1001400 0 180 $X=974020 $Y=995980
X2053 5783 5328 5719 2 1 5776 QDFFRBN $T=975880 1011480 1 0 $X=975880 $Y=1006060
X2054 5766 973 5790 2 1 5778 QDFFRBN $T=988280 951000 0 180 $X=976500 $Y=945580
X2055 5789 973 5697 2 1 1079 QDFFRBN $T=977740 961080 0 0 $X=977740 $Y=960700
X2056 5781 5328 5717 2 1 5734 QDFFRBN $T=989520 1041720 0 180 $X=977740 $Y=1036300
X2057 5806 5328 5743 2 1 1051 QDFFRBN $T=990760 1041720 1 180 $X=978980 $Y=1041340
X2058 5793 973 5732 2 1 1081 QDFFRBN $T=979600 951000 0 0 $X=979600 $Y=950620
X2059 5832 5328 5743 2 1 5791 QDFFRBN $T=991380 1031640 0 180 $X=979600 $Y=1026220
X2060 5799 946 5763 2 1 5841 QDFFRBN $T=980220 1061880 0 0 $X=980220 $Y=1061500
X2061 5800 946 1076 2 1 5842 QDFFRBN $T=980220 1082040 1 0 $X=980220 $Y=1076620
X2062 5803 973 1078 2 1 5824 QDFFRBN $T=980840 910680 0 0 $X=980840 $Y=910300
X2063 5812 5328 5847 2 1 1085 QDFFRBN $T=983940 1051800 1 0 $X=983940 $Y=1046380
X2064 5859 946 5763 2 1 5808 QDFFRBN $T=995720 1061880 0 180 $X=983940 $Y=1056460
X2065 5814 5328 5719 2 1 5833 QDFFRBN $T=984560 1001400 0 0 $X=984560 $Y=1001020
X2066 5815 5328 5804 2 1 5813 QDFFRBN $T=984560 1011480 0 0 $X=984560 $Y=1011100
X2067 5825 5328 5854 2 1 5823 QDFFRBN $T=987040 981240 1 0 $X=987040 $Y=975820
X2068 5826 973 1078 2 1 5885 QDFFRBN $T=987660 920760 1 0 $X=987660 $Y=915340
X2069 5831 973 1078 2 1 5889 QDFFRBN $T=989520 910680 1 0 $X=989520 $Y=905260
X2070 5838 973 5872 2 1 5865 QDFFRBN $T=990140 951000 1 0 $X=990140 $Y=945580
X2071 5834 5328 5854 2 1 5893 QDFFRBN $T=990140 991320 1 0 $X=990140 $Y=985900
X2072 5844 5328 5719 2 1 5890 QDFFRBN $T=991380 1001400 1 0 $X=991380 $Y=995980
X2073 5882 5328 5847 2 1 5820 QDFFRBN $T=1003160 1041720 0 180 $X=991380 $Y=1036300
X2074 5848 5328 5872 2 1 5855 QDFFRBN $T=992000 971160 1 0 $X=992000 $Y=965740
X2075 5850 973 5872 2 1 5874 QDFFRBN $T=992620 951000 0 0 $X=992620 $Y=950620
X2076 5863 946 5910 2 1 5924 QDFFRBN $T=995100 1051800 0 0 $X=995100 $Y=1051420
X2077 5878 973 5765 2 1 5819 QDFFRBN $T=998200 920760 0 0 $X=998200 $Y=920380
X2078 5880 5328 5804 2 1 5932 QDFFRBN $T=998200 1011480 0 0 $X=998200 $Y=1011100
X2079 5954 1115 5765 2 1 5886 QDFFRBN $T=1011840 930840 0 180 $X=1000060 $Y=925420
X2080 5912 5328 5854 2 1 5836 QDFFRBN $T=1003160 981240 0 0 $X=1003160 $Y=980860
X2081 5914 973 5872 2 1 5982 QDFFRBN $T=1003780 951000 1 0 $X=1003780 $Y=945580
X2082 5926 973 5872 2 1 1133 QDFFRBN $T=1004400 961080 0 0 $X=1004400 $Y=960700
X2083 5927 5328 5975 2 1 5985 QDFFRBN $T=1005020 1001400 0 0 $X=1005020 $Y=1001020
X2084 5966 1115 1086 2 1 1106 QDFFRBN $T=1017420 900600 1 180 $X=1005640 $Y=900220
X2085 5908 973 5872 2 1 5929 QDFFRBN $T=1006260 971160 1 0 $X=1006260 $Y=965740
X2086 5935 5328 5854 2 1 1131 QDFFRBN $T=1006260 991320 1 0 $X=1006260 $Y=985900
X2087 5950 5328 5975 2 1 5974 QDFFRBN $T=1009360 1031640 1 0 $X=1009360 $Y=1026220
X2088 5951 946 5910 2 1 5965 QDFFRBN $T=1009360 1051800 0 0 $X=1009360 $Y=1051420
X2089 5979 5328 5975 2 1 5963 QDFFRBN $T=1023000 1031640 1 180 $X=1011220 $Y=1031260
X2090 5967 1115 6018 2 1 5987 QDFFRBN $T=1011840 920760 0 0 $X=1011840 $Y=920380
X2091 5970 5328 6020 2 1 5960 QDFFRBN $T=1011840 1011480 0 0 $X=1011840 $Y=1011100
X2092 5981 1115 5938 2 1 1143 QDFFRBN $T=1014320 930840 1 0 $X=1014320 $Y=925420
X2093 6047 6041 5854 2 1 5996 QDFFRBN $T=1028580 981240 1 180 $X=1016800 $Y=980860
X2094 5989 1149 1135 2 1 1098 QDFFRBN $T=1028580 1082040 1 180 $X=1016800 $Y=1081660
X2095 1138 1115 6018 2 1 1152 QDFFRBN $T=1018660 900600 0 0 $X=1018660 $Y=900220
X2096 6056 1115 6018 2 1 6012 QDFFRBN $T=1031060 920760 0 180 $X=1019280 $Y=915340
X2097 6048 6041 6029 2 1 5957 QDFFRBN $T=1031680 961080 1 180 $X=1019900 $Y=960700
X2098 6042 6041 6029 2 1 6019 QDFFRBN $T=1031680 971160 1 180 $X=1019900 $Y=970780
X2099 6021 5328 6020 2 1 1144 QDFFRBN $T=1019900 1001400 0 0 $X=1019900 $Y=1001020
X2100 6068 1149 1118 2 1 6022 QDFFRBN $T=1032300 1061880 0 180 $X=1020520 $Y=1056460
X2101 6077 1115 5938 2 1 1141 QDFFRBN $T=1034160 930840 1 180 $X=1022380 $Y=930460
X2102 6067 6041 6029 2 1 6025 QDFFRBN $T=1034160 951000 1 180 $X=1022380 $Y=950620
X2103 6066 6041 5975 2 1 6032 QDFFRBN $T=1035400 1021560 1 180 $X=1023620 $Y=1021180
X2104 6037 6041 6020 2 1 6036 QDFFRBN $T=1024240 1031640 1 0 $X=1024240 $Y=1026220
X2105 6090 6041 5975 2 1 6017 QDFFRBN $T=1036640 1031640 1 180 $X=1024860 $Y=1031260
X2106 6043 6041 5975 2 1 6040 QDFFRBN $T=1037260 1011480 1 180 $X=1025480 $Y=1011100
X2107 6103 1115 5938 2 1 5990 QDFFRBN $T=1038500 930840 0 180 $X=1026720 $Y=925420
X2108 6049 946 6093 2 1 6098 QDFFRBN $T=1027340 1071960 1 0 $X=1027340 $Y=1066540
X2109 6065 6041 6020 2 1 6023 QDFFRBN $T=1039740 991320 1 180 $X=1027960 $Y=990940
X2110 6062 1149 6093 2 1 5980 QDFFRBN $T=1029200 1051800 0 0 $X=1029200 $Y=1051420
X2111 1155 1149 1118 2 1 1167 QDFFRBN $T=1030440 1082040 0 0 $X=1030440 $Y=1081660
X2112 6053 1115 6018 2 1 1128 QDFFRBN $T=1043460 900600 1 180 $X=1031680 $Y=900220
X2113 6085 6041 6126 2 1 6009 QDFFRBN $T=1033540 981240 1 0 $X=1033540 $Y=975820
X2114 6094 6041 6029 2 1 1178 QDFFRBN $T=1035400 971160 0 0 $X=1035400 $Y=970780
X2115 6104 6041 6144 2 1 6132 QDFFRBN $T=1036640 1021560 1 0 $X=1036640 $Y=1016140
X2116 6107 1115 6146 2 1 6074 QDFFRBN $T=1037260 940920 0 0 $X=1037260 $Y=940540
X2117 6115 1115 5938 2 1 6165 QDFFRBN $T=1039120 930840 1 0 $X=1039120 $Y=925420
X2118 6121 1115 5938 2 1 6139 QDFFRBN $T=1040360 930840 0 0 $X=1040360 $Y=930460
X2119 6172 1149 1118 2 1 6128 QDFFRBN $T=1054000 1071960 0 180 $X=1042220 $Y=1066540
X2120 6177 1115 1161 2 1 6135 QDFFRBN $T=1054620 910680 0 180 $X=1042840 $Y=905260
X2121 6129 1115 6167 2 1 1158 QDFFRBN $T=1042840 920760 1 0 $X=1042840 $Y=915340
X2122 6182 1149 5910 2 1 6134 QDFFRBN $T=1054620 1051800 1 180 $X=1042840 $Y=1051420
X2123 6114 6041 6144 2 1 6138 QDFFRBN $T=1056480 1001400 1 180 $X=1044700 $Y=1001020
X2124 6156 1149 6187 2 1 6073 QDFFRBN $T=1046560 1041720 0 0 $X=1046560 $Y=1041340
X2125 6160 6041 6162 2 1 6203 QDFFRBN $T=1047800 961080 1 0 $X=1047800 $Y=955660
X2126 6131 6041 6126 2 1 6143 QDFFRBN $T=1059580 1001400 0 180 $X=1047800 $Y=995980
X2127 6163 1149 6194 2 1 6124 QDFFRBN $T=1047800 1041720 1 0 $X=1047800 $Y=1036300
X2128 6147 1149 6187 2 1 6079 QDFFRBN $T=1049040 1051800 1 0 $X=1049040 $Y=1046380
X2129 6216 1115 1161 2 1 1184 QDFFRBN $T=1062680 910680 1 180 $X=1050900 $Y=910300
X2130 6166 6041 6144 2 1 1172 QDFFRBN $T=1062680 1011480 1 180 $X=1050900 $Y=1011100
X2131 1203 1149 6093 2 1 1185 QDFFRBN $T=1062680 1082040 0 180 $X=1050900 $Y=1076620
X2132 6154 6041 6144 2 1 1164 QDFFRBN $T=1063300 1021560 0 180 $X=1051520 $Y=1016140
X2133 6178 6041 6126 2 1 6210 QDFFRBN $T=1052760 991320 0 0 $X=1052760 $Y=990940
X2134 6179 1149 1198 2 1 1174 QDFFRBN $T=1052760 1071960 0 0 $X=1052760 $Y=1071580
X2135 6195 1115 6167 2 1 6237 QDFFRBN $T=1055860 910680 1 0 $X=1055860 $Y=905260
X2136 6207 6041 6259 2 1 6248 QDFFRBN $T=1058960 981240 0 0 $X=1058960 $Y=980860
X2137 6208 6041 6126 2 1 6225 QDFFRBN $T=1058960 1001400 0 0 $X=1058960 $Y=1001020
X2138 6263 6041 6187 2 1 6209 QDFFRBN $T=1071360 1031640 0 180 $X=1059580 $Y=1026220
X2139 6273 1149 1198 2 1 6221 QDFFRBN $T=1072600 1041720 1 180 $X=1060820 $Y=1041340
X2140 6222 6041 6194 2 1 6281 QDFFRBN $T=1061440 1021560 0 0 $X=1061440 $Y=1021180
X2141 6278 6041 6162 2 1 6224 QDFFRBN $T=1073840 971160 0 180 $X=1062060 $Y=965740
X2142 6215 1149 6236 2 1 1206 QDFFRBN $T=1075700 1051800 1 180 $X=1063920 $Y=1051420
X2143 6242 1149 1198 2 1 6267 QDFFRBN $T=1063920 1082040 1 0 $X=1063920 $Y=1076620
X2144 6247 1149 6236 2 1 6293 QDFFRBN $T=1064540 1071960 0 0 $X=1064540 $Y=1071580
X2145 6229 1115 6167 2 1 1202 QDFFRBN $T=1076940 930840 0 180 $X=1065160 $Y=925420
X2146 6286 6041 6146 2 1 6251 QDFFRBN $T=1077560 940920 1 180 $X=1065780 $Y=940540
X2147 6258 6041 6259 2 1 1219 QDFFRBN $T=1066400 991320 0 0 $X=1066400 $Y=990940
X2148 6252 1115 6146 2 1 6213 QDFFRBN $T=1078800 930840 1 180 $X=1067020 $Y=930460
X2149 6301 6041 6259 2 1 6260 QDFFRBN $T=1078800 991320 0 180 $X=1067020 $Y=985900
X2150 6270 6041 6259 2 1 1226 QDFFRBN $T=1068880 1001400 1 0 $X=1068880 $Y=995980
X2151 6272 6041 6194 2 1 6243 QDFFRBN $T=1073220 1021560 0 0 $X=1073220 $Y=1021180
X2152 6264 1149 6236 2 1 6284 QDFFRBN $T=1073220 1041720 1 0 $X=1073220 $Y=1036300
X2153 6276 1149 6236 2 1 6220 QDFFRBN $T=1073840 1041720 0 0 $X=1073840 $Y=1041340
X2154 6296 1115 6332 2 1 6350 QDFFRBN $T=1076320 920760 0 0 $X=1076320 $Y=920380
X2155 6302 1149 6333 2 1 6322 QDFFRBN $T=1076940 1051800 0 0 $X=1076940 $Y=1051420
X2156 1220 1115 1212 2 1 1201 QDFFRBN $T=1077560 910680 1 0 $X=1077560 $Y=905260
X2157 6310 6041 6346 2 1 6291 QDFFRBN $T=1079420 1011480 0 0 $X=1079420 $Y=1011100
X2158 6314 6041 6336 2 1 6351 QDFFRBN $T=1080040 981240 0 0 $X=1080040 $Y=980860
X2159 6318 6041 6336 2 1 6294 QDFFRBN $T=1080660 971160 0 0 $X=1080660 $Y=970780
X2160 6319 6041 6346 2 1 6376 QDFFRBN $T=1080660 1011480 1 0 $X=1080660 $Y=1006060
X2161 6326 6041 6336 2 1 6298 QDFFRBN $T=1081900 961080 0 0 $X=1081900 $Y=960700
X2162 6372 6041 6336 2 1 6328 QDFFRBN $T=1093680 991320 1 180 $X=1081900 $Y=990940
X2163 6327 6041 6336 2 1 1213 QDFFRBN $T=1095540 971160 0 180 $X=1083760 $Y=965740
X2164 6337 1149 6194 2 1 6373 QDFFRBN $T=1085000 1021560 0 0 $X=1085000 $Y=1021180
X2165 6394 1149 6333 2 1 1231 QDFFRBN $T=1098020 1051800 0 180 $X=1086240 $Y=1046380
X2166 6353 1149 6194 2 1 6360 QDFFRBN $T=1087480 1041720 0 0 $X=1087480 $Y=1041340
X2167 6355 1115 1212 2 1 1254 QDFFRBN $T=1088100 920760 1 0 $X=1088100 $Y=915340
X2168 6356 6041 6398 2 1 6371 QDFFRBN $T=1088100 981240 1 0 $X=1088100 $Y=975820
X2169 6358 1115 1212 2 1 1253 QDFFRBN $T=1088720 910680 0 0 $X=1088720 $Y=910300
X2170 6377 1115 6332 2 1 6320 QDFFRBN $T=1101740 920760 1 180 $X=1089960 $Y=920380
X2171 6417 1149 6333 2 1 1237 QDFFRBN $T=1102360 1051800 1 180 $X=1090580 $Y=1051420
X2172 6374 6041 6312 2 1 6343 QDFFRBN $T=1102980 940920 0 180 $X=1091200 $Y=935500
X2173 6362 6041 6312 2 1 6344 QDFFRBN $T=1093060 940920 0 0 $X=1093060 $Y=940540
X2174 6392 1149 1250 2 1 6436 QDFFRBN $T=1094920 1071960 0 0 $X=1094920 $Y=1071580
X2175 6445 1149 1250 2 1 6395 QDFFRBN $T=1107320 1082040 1 180 $X=1095540 $Y=1081660
X2176 6410 6041 6346 2 1 6405 QDFFRBN $T=1098020 1011480 1 0 $X=1098020 $Y=1006060
X2177 6428 1149 6450 2 1 6331 QDFFRBN $T=1101120 1041720 1 0 $X=1101120 $Y=1036300
X2178 6458 1149 6333 2 1 6418 QDFFRBN $T=1112900 1041720 1 180 $X=1101120 $Y=1041340
X2179 6489 1115 6167 2 1 6433 QDFFRBN $T=1114760 910680 0 180 $X=1102980 $Y=905260
X2180 6438 1115 6332 2 1 6457 QDFFRBN $T=1103600 920760 0 0 $X=1103600 $Y=920380
X2181 6455 6041 6312 2 1 6413 QDFFRBN $T=1115380 940920 0 180 $X=1103600 $Y=935500
X2182 6429 6041 6398 2 1 1262 QDFFRBN $T=1115380 971160 1 180 $X=1103600 $Y=970780
X2183 6481 6041 6398 2 1 6414 QDFFRBN $T=1115380 981240 1 180 $X=1103600 $Y=980860
X2184 6465 1149 6450 2 1 6427 QDFFRBN $T=1115380 1021560 1 180 $X=1103600 $Y=1021180
X2185 6495 6041 6398 2 1 6439 QDFFRBN $T=1116000 961080 0 180 $X=1104220 $Y=955660
X2186 6496 6041 6398 2 1 6452 QDFFRBN $T=1119100 961080 1 180 $X=1107320 $Y=960700
X2187 6462 6041 6346 2 1 6453 QDFFRBN $T=1108560 1001400 0 0 $X=1108560 $Y=1001020
X2188 6521 6041 6477 2 1 6461 QDFFRBN $T=1123440 940920 1 180 $X=1111660 $Y=940540
X2189 6515 1115 1214 2 1 1275 QDFFRBN $T=1128400 910680 0 180 $X=1116620 $Y=905260
X2190 6527 6041 6332 2 1 6485 QDFFRBN $T=1128400 920760 0 180 $X=1116620 $Y=915340
X2191 6497 6041 1282 2 1 6430 QDFFRBN $T=1128400 930840 0 180 $X=1116620 $Y=925420
X2192 6528 6041 6477 2 1 6505 QDFFRBN $T=1128400 940920 0 180 $X=1116620 $Y=935500
X2193 6507 6041 6477 2 1 6500 QDFFRBN $T=1128400 981240 1 180 $X=1116620 $Y=980860
X2194 6523 6041 6477 2 1 6506 QDFFRBN $T=1128400 991320 0 180 $X=1116620 $Y=985900
X2195 6529 6041 6346 2 1 6501 QDFFRBN $T=1128400 1001400 0 180 $X=1116620 $Y=995980
X2196 6508 6041 6450 2 1 6421 QDFFRBN $T=1128400 1011480 0 180 $X=1116620 $Y=1006060
X2197 6524 1149 6450 2 1 6471 QDFFRBN $T=1128400 1021560 1 180 $X=1116620 $Y=1021180
X2198 6504 1149 1250 2 1 6460 QDFFRBN $T=1128400 1071960 1 180 $X=1116620 $Y=1071580
X2199 6494 1149 1250 2 1 6463 QDFFRBN $T=1128400 1082040 0 180 $X=1116620 $Y=1076620
X2200 6530 6041 6477 2 1 6509 QDFFRBN $T=1129020 961080 0 180 $X=1117240 $Y=955660
X2201 6514 1149 6512 2 1 6487 QDFFRBN $T=1129020 1041720 1 180 $X=1117240 $Y=1041340
X2202 6498 1149 6512 2 1 6469 QDFFRBN $T=1129020 1071960 0 180 $X=1117240 $Y=1066540
X2203 6531 6041 6477 2 1 6513 QDFFRBN $T=1129640 971160 0 180 $X=1117860 $Y=965740
X2204 6511 1149 6450 2 1 6482 QDFFRBN $T=1129640 1031640 1 180 $X=1117860 $Y=1031260
X2205 6503 1149 6512 2 1 6448 QDFFRBN $T=1129640 1051800 1 180 $X=1117860 $Y=1051420
X2206 2243 1 2 2267 2274 2307 1299 ICV_4 $T=361460 1031640 0 0 $X=361460 $Y=1031260
X2207 2292 1 2 2325 2330 2360 1299 ICV_4 $T=368900 1071960 0 0 $X=368900 $Y=1071580
X2208 2313 1 2 2344 2349 2370 1299 ICV_4 $T=371380 1031640 0 0 $X=371380 $Y=1031260
X2209 2355 1 2 2384 2381 2416 1299 ICV_4 $T=378820 1071960 0 0 $X=378820 $Y=1071580
X2210 2390 1 2 2414 2406 2442 1299 ICV_4 $T=383160 1031640 1 0 $X=383160 $Y=1026220
X2211 2374 1 2 2391 2356 2415 1299 ICV_4 $T=383780 1051800 0 0 $X=383780 $Y=1051420
X2212 2457 1 2 2490 2493 2519 1299 ICV_4 $T=395560 1051800 0 0 $X=395560 $Y=1051420
X2213 2501 1 2 2533 2498 2573 1299 ICV_4 $T=402380 981240 0 0 $X=402380 $Y=980860
X2214 2597 1 2 2625 2631 2653 1299 ICV_4 $T=416020 910680 1 0 $X=416020 $Y=905260
X2215 2660 1 2 2686 2687 2712 1299 ICV_4 $T=425940 910680 1 0 $X=425940 $Y=905260
X2216 2674 1 2 2698 2703 2731 1299 ICV_4 $T=428420 951000 1 0 $X=428420 $Y=945580
X2217 2668 1 2 2663 2709 2736 1299 ICV_4 $T=429660 1051800 1 0 $X=429660 $Y=1046380
X2218 2717 1 2 261 2742 2765 1299 ICV_4 $T=435860 910680 1 0 $X=435860 $Y=905260
X2219 2817 1 2 2792 2833 2837 1299 ICV_4 $T=453840 961080 0 0 $X=453840 $Y=960700
X2220 2869 1 2 2873 298 2905 1299 ICV_4 $T=463760 1071960 1 0 $X=463760 $Y=1066540
X2221 2880 1 2 2871 2907 2857 1299 ICV_4 $T=465620 1021560 1 0 $X=465620 $Y=1016140
X2222 2963 1 2 2988 2985 3011 1299 ICV_4 $T=480500 1021560 1 0 $X=480500 $Y=1016140
X2223 2973 1 2 2983 2999 3028 1299 ICV_4 $T=482360 1061880 1 0 $X=482360 $Y=1056460
X2224 2962 1 2 2938 2974 3006 1299 ICV_4 $T=484220 961080 1 0 $X=484220 $Y=955660
X2225 2996 1 2 3017 3026 3016 1299 ICV_4 $T=490420 1021560 1 0 $X=490420 $Y=1016140
X2226 3018 1 2 3045 2959 3072 1299 ICV_4 $T=491040 961080 0 0 $X=491040 $Y=960700
X2227 3020 1 2 3051 3117 3105 1299 ICV_4 $T=504060 991320 1 0 $X=504060 $Y=985900
X2228 328 1 2 3110 3112 3140 1299 ICV_4 $T=506540 920760 1 0 $X=506540 $Y=915340
X2229 3199 1 2 3198 3218 3241 1299 ICV_4 $T=523900 991320 1 0 $X=523900 $Y=985900
X2230 3151 1 2 3200 2989 3001 1299 ICV_4 $T=523900 1011480 0 0 $X=523900 $Y=1011100
X2231 370 1 2 3263 3275 3298 1299 ICV_4 $T=533820 920760 1 0 $X=533820 $Y=915340
X2232 3250 1 2 3249 3174 3225 1299 ICV_4 $T=534440 1082040 1 0 $X=534440 $Y=1076620
X2233 3189 1 2 3215 3284 3254 1299 ICV_4 $T=535680 1021560 1 0 $X=535680 $Y=1016140
X2234 3315 1 2 3337 3339 3347 1299 ICV_4 $T=544980 971160 1 0 $X=544980 $Y=965740
X2235 3126 1 2 3152 3344 3332 1299 ICV_4 $T=545600 1021560 1 0 $X=545600 $Y=1016140
X2236 3260 1 2 3296 3357 3375 1299 ICV_4 $T=546840 1061880 0 0 $X=546840 $Y=1061500
X2237 3322 1 2 3349 410 3361 1299 ICV_4 $T=546840 1082040 1 0 $X=546840 $Y=1076620
X2238 3355 1 2 3382 3408 3425 1299 ICV_4 $T=556140 981240 1 0 $X=556140 $Y=975820
X2239 3435 1 2 3451 3462 3485 1299 ICV_4 $T=566680 920760 0 0 $X=566680 $Y=920380
X2240 3371 1 2 3352 3235 3265 1299 ICV_4 $T=568540 1041720 1 0 $X=568540 $Y=1036300
X2241 3448 1 2 3474 3412 3467 1299 ICV_4 $T=573500 1071960 1 0 $X=573500 $Y=1066540
X2242 3487 1 2 3505 3510 3538 1299 ICV_4 $T=577220 1011480 1 0 $X=577220 $Y=1006060
X2243 448 1 2 3543 3527 3536 1299 ICV_4 $T=585280 1071960 0 0 $X=585280 $Y=1071580
X2244 3550 1 2 3568 3569 3590 1299 ICV_4 $T=590240 1011480 1 0 $X=590240 $Y=1006060
X2245 3466 1 2 3402 3573 3594 1299 ICV_4 $T=590860 930840 0 0 $X=590860 $Y=930460
X2246 3546 1 2 3562 3577 3595 1299 ICV_4 $T=590860 961080 0 0 $X=590860 $Y=960700
X2247 3563 1 2 3583 3588 3608 1299 ICV_4 $T=593960 1021560 0 0 $X=593960 $Y=1021180
X2248 3570 1 2 3591 3596 3614 1299 ICV_4 $T=595200 1051800 1 0 $X=595200 $Y=1046380
X2249 3571 1 2 3600 3602 3624 1299 ICV_4 $T=596440 1071960 0 0 $X=596440 $Y=1071580
X2250 491 1 2 497 3621 3649 1299 ICV_4 $T=601400 900600 0 0 $X=601400 $Y=900220
X2251 3609 1 2 3637 3643 3663 1299 ICV_4 $T=603880 940920 1 0 $X=603880 $Y=935500
X2252 3603 1 2 3645 3589 3665 1299 ICV_4 $T=612560 930840 0 0 $X=612560 $Y=930460
X2253 3612 1 2 3683 3744 3767 1299 ICV_4 $T=619380 1061880 1 0 $X=619380 $Y=1056460
X2254 3728 1 2 3740 3691 3750 1299 ICV_4 $T=622480 930840 0 0 $X=622480 $Y=930460
X2255 3733 1 2 3762 3766 3789 1299 ICV_4 $T=623720 1001400 0 0 $X=623720 $Y=1001020
X2256 3820 1 2 3833 3855 3871 1299 ICV_4 $T=643560 1071960 0 0 $X=643560 $Y=1071580
X2257 3899 1 2 3889 3908 3912 1299 ICV_4 $T=658440 1051800 0 0 $X=658440 $Y=1051420
X2258 3902 1 2 3893 3945 3979 1299 ICV_4 $T=659680 930840 0 0 $X=659680 $Y=930460
X2259 3949 1 2 3985 3992 4013 1299 ICV_4 $T=665260 991320 0 0 $X=665260 $Y=990940
X2260 3934 1 2 3952 3978 3956 1299 ICV_4 $T=665260 1031640 1 0 $X=665260 $Y=1026220
X2261 3954 1 2 3988 3993 4017 1299 ICV_4 $T=665880 951000 0 0 $X=665880 $Y=950620
X2262 4012 1 2 4039 4046 4071 1299 ICV_4 $T=674560 981240 0 0 $X=674560 $Y=980860
X2263 4052 1 2 4084 638 4112 1299 ICV_4 $T=681380 1061880 1 0 $X=681380 $Y=1056460
X2264 4043 1 2 4077 4063 4096 1299 ICV_4 $T=684480 981240 0 0 $X=684480 $Y=980860
X2265 4127 1 2 4177 4198 4205 1299 ICV_4 $T=699980 981240 0 0 $X=699980 $Y=980860
X2266 4195 1 2 4220 4178 4229 1299 ICV_4 $T=705560 1041720 0 0 $X=705560 $Y=1041340
X2267 4233 1 2 4262 4270 4295 1299 ICV_4 $T=714860 930840 0 0 $X=714860 $Y=930460
X2268 4223 1 2 4245 4252 4228 1299 ICV_4 $T=714860 961080 1 0 $X=714860 $Y=955660
X2269 4285 1 2 4280 4277 4318 1299 ICV_4 $T=722920 1041720 0 0 $X=722920 $Y=1041340
X2270 4370 1 2 4369 4333 4347 1299 ICV_4 $T=734080 1041720 0 0 $X=734080 $Y=1041340
X2271 4301 1 2 4358 4140 4202 1299 ICV_4 $T=736560 930840 0 0 $X=736560 $Y=930460
X2272 4337 1 2 4398 4377 4437 1299 ICV_4 $T=744000 1041720 0 0 $X=744000 $Y=1041340
X2273 4394 1 2 4396 4345 4392 1299 ICV_4 $T=749580 940920 1 0 $X=749580 $Y=935500
X2274 4456 1 2 4481 4487 4509 1299 ICV_4 $T=752680 1011480 1 0 $X=752680 $Y=1006060
X2275 4483 1 2 4507 4512 4519 1299 ICV_4 $T=757020 1071960 0 0 $X=757020 $Y=1071580
X2276 4676 1 2 4701 4713 4745 1299 ICV_4 $T=788020 951000 1 0 $X=788020 $Y=945580
X2277 4750 1 2 4777 4783 4812 1299 ICV_4 $T=797940 951000 1 0 $X=797940 $Y=945580
X2278 4760 1 2 4785 4772 4834 1299 ICV_4 $T=799800 910680 1 0 $X=799800 $Y=905260
X2279 4323 1 2 4314 4800 4801 1299 ICV_4 $T=800420 1051800 0 0 $X=800420 $Y=1051420
X2280 4847 1 2 4787 4786 4811 1299 ICV_4 $T=812200 1061880 1 0 $X=812200 $Y=1056460
X2281 4733 1 2 4796 4863 4864 1299 ICV_4 $T=819020 1011480 1 0 $X=819020 $Y=1006060
X2282 4822 1 2 4804 4689 4814 1299 ICV_4 $T=819020 1041720 0 0 $X=819020 $Y=1041340
X2283 4915 1 2 4919 4769 4791 1299 ICV_4 $T=825840 1061880 0 0 $X=825840 $Y=1061500
X2284 4916 1 2 4950 4953 4978 1299 ICV_4 $T=827080 1051800 1 0 $X=827080 $Y=1046380
X2285 4947 1 2 4956 4976 4981 1299 ICV_4 $T=831420 1011480 0 0 $X=831420 $Y=1011100
X2286 5005 1 2 5023 5036 5035 1299 ICV_4 $T=841340 1051800 0 0 $X=841340 $Y=1051420
X2287 4941 1 2 5017 5015 5053 1299 ICV_4 $T=846300 981240 1 0 $X=846300 $Y=975820
X2288 5123 1 2 5170 5154 5194 1299 ICV_4 $T=865520 1061880 1 0 $X=865520 $Y=1056460
X2289 5171 1 2 5197 5202 5211 1299 ICV_4 $T=869240 971160 1 0 $X=869240 $Y=965740
X2290 5175 1 2 5201 5209 5208 1299 ICV_4 $T=869860 930840 0 0 $X=869860 $Y=930460
X2291 910 1 2 913 5136 5219 1299 ICV_4 $T=872340 1082040 1 0 $X=872340 $Y=1076620
X2292 5199 1 2 5230 5235 5234 1299 ICV_4 $T=874200 1051800 0 0 $X=874200 $Y=1051420
X2293 5253 1 2 5238 5290 5232 1299 ICV_4 $T=882260 1082040 1 0 $X=882260 $Y=1076620
X2294 5243 1 2 5285 5193 5217 1299 ICV_4 $T=884120 1021560 1 0 $X=884120 $Y=1016140
X2295 5203 1 2 5260 5259 5317 1299 ICV_4 $T=887220 991320 0 0 $X=887220 $Y=990940
X2296 5305 1 2 5329 5311 5337 1299 ICV_4 $T=889080 900600 0 0 $X=889080 $Y=900220
X2297 5299 1 2 5339 5345 5371 1299 ICV_4 $T=891560 940920 0 0 $X=891560 $Y=940540
X2298 5375 1 2 5392 5397 5396 1299 ICV_4 $T=901480 981240 1 0 $X=901480 $Y=975820
X2299 5367 1 2 5376 5330 5295 1299 ICV_4 $T=901480 1001400 0 0 $X=901480 $Y=1001020
X2300 964 1 2 968 5380 5390 1299 ICV_4 $T=908920 910680 1 0 $X=908920 $Y=905260
X2301 5137 1 2 5127 5091 5113 1299 ICV_4 $T=908920 961080 1 0 $X=908920 $Y=955660
X2302 5407 1 2 5428 5424 5448 1299 ICV_4 $T=910160 1061880 1 0 $X=910160 $Y=1056460
X2303 5413 1 2 5389 5417 5426 1299 ICV_4 $T=913260 1001400 1 0 $X=913260 $Y=995980
X2304 5383 1 2 5425 5447 5480 1299 ICV_4 $T=914500 1031640 0 0 $X=914500 $Y=1031260
X2305 5491 1 2 5506 5512 5518 1299 ICV_4 $T=925040 930840 1 0 $X=925040 $Y=925420
X2306 992 1 2 1003 5483 5492 1299 ICV_4 $T=926900 1082040 1 0 $X=926900 $Y=1076620
X2307 5507 1 2 5536 5539 5538 1299 ICV_4 $T=929380 1001400 1 0 $X=929380 $Y=995980
X2308 5573 1 2 5542 5602 5604 1299 ICV_4 $T=939300 1001400 1 0 $X=939300 $Y=995980
X2309 5582 1 2 5597 5520 5554 1299 ICV_4 $T=943640 961080 0 0 $X=943640 $Y=960700
X2310 5612 1 2 5608 1030 1037 1299 ICV_4 $T=947360 910680 0 0 $X=947360 $Y=910300
X2311 5623 1 2 5640 5639 5659 1299 ICV_4 $T=947980 1061880 1 0 $X=947980 $Y=1056460
X2312 5616 1 2 5664 1055 1061 1299 ICV_4 $T=960380 900600 0 0 $X=960380 $Y=900220
X2313 5699 1 2 5723 5730 5731 1299 ICV_4 $T=960380 1061880 1 0 $X=960380 $Y=1056460
X2314 1054 1 2 1064 1066 1069 1299 ICV_4 $T=965340 1082040 0 0 $X=965340 $Y=1081660
X2315 5684 1 2 5733 5722 5759 1299 ICV_4 $T=965960 1031640 0 0 $X=965960 $Y=1031260
X2316 5736 1 2 1071 5741 5774 1299 ICV_4 $T=972160 910680 1 0 $X=972160 $Y=905260
X2317 5767 1 2 5784 5768 5801 1299 ICV_4 $T=975880 971160 0 0 $X=975880 $Y=970780
X2318 5725 1 2 5782 5702 5739 1299 ICV_4 $T=975880 1082040 0 0 $X=975880 $Y=1081660
X2319 5805 1 2 5818 5820 5845 1299 ICV_4 $T=981460 1031640 0 0 $X=981460 $Y=1031260
X2320 5813 1 2 5830 5833 5837 1299 ICV_4 $T=985180 1021560 1 0 $X=985180 $Y=1016140
X2321 5855 1 2 5869 5874 5873 1299 ICV_4 $T=993240 961080 0 0 $X=993240 $Y=960700
X2322 5893 1 2 5875 5890 5876 1299 ICV_4 $T=1003780 991320 0 0 $X=1003780 $Y=990940
X2323 5808 1 2 5895 5934 5945 1299 ICV_4 $T=1016800 1082040 1 0 $X=1016800 $Y=1076620
X2324 6009 1 2 6030 6019 6033 1299 ICV_4 $T=1018660 971160 1 0 $X=1018660 $Y=965740
X2325 5963 1 2 5953 6017 6069 1299 ICV_4 $T=1022380 1041720 1 0 $X=1022380 $Y=1036300
X2326 6012 1 2 6038 5681 5716 1299 ICV_4 $T=1024860 910680 1 0 $X=1024860 $Y=905260
X2327 6098 1 2 6117 6128 6152 1299 ICV_4 $T=1036640 1082040 1 0 $X=1036640 $Y=1076620
X2328 1167 1 2 1175 1177 1186 1299 ICV_4 $T=1042220 1082040 0 0 $X=1042220 $Y=1081660
X2329 6221 1 2 6250 6267 6266 1299 ICV_4 $T=1062680 1082040 0 0 $X=1062680 $Y=1081660
X2330 6251 1 2 6275 6203 6180 1299 ICV_4 $T=1065780 951000 0 0 $X=1065780 $Y=950620
X2331 6257 1 2 6283 6293 6282 1299 ICV_4 $T=1070740 1061880 1 0 $X=1070740 $Y=1056460
X2332 6260 1 2 6289 6294 6306 1299 ICV_4 $T=1078800 991320 1 0 $X=1078800 $Y=985900
X2333 6320 1 2 6341 6344 6345 1299 ICV_4 $T=1081280 940920 1 0 $X=1081280 $Y=935500
X2334 6298 1 2 6308 6351 6335 1299 ICV_4 $T=1082520 961080 1 0 $X=1082520 $Y=955660
X2335 6331 1 2 6357 6360 6385 1299 ICV_4 $T=1084380 1031640 0 0 $X=1084380 $Y=1031260
X2336 6339 1 2 6364 6386 6387 1299 ICV_4 $T=1089340 1061880 1 0 $X=1089340 $Y=1056460
X2337 6381 1 2 6383 6248 6219 1299 ICV_4 $T=1094300 961080 1 0 $X=1094300 $Y=955660
X2338 1261 1 2 1271 6457 6464 1299 ICV_4 $T=1103600 910680 0 0 $X=1103600 $Y=910300
X2339 6485 1 2 6516 1283 1285 1299 ICV_4 $T=1115380 920760 0 0 $X=1115380 $Y=920380
X2340 6418 1 2 6443 6311 6347 1299 ICV_4 $T=1116620 1051800 1 0 $X=1116620 $Y=1046380
X2341 6471 1 2 6518 6281 6256 1299 ICV_4 $T=1118480 1021560 1 0 $X=1118480 $Y=1016140
X2342 6487 1 2 6493 6427 6444 1299 ICV_4 $T=1118480 1041720 1 0 $X=1118480 $Y=1036300
X2343 6436 1 2 6459 6469 6476 1299 ICV_4 $T=1118480 1061880 0 0 $X=1118480 $Y=1061500
X2344 6501 1 2 6522 6513 6526 1299 ICV_4 $T=1119720 981240 1 0 $X=1119720 $Y=975820
X2345 2384 2385 2 1 2278 193 MUX2 $T=383160 1061880 1 180 $X=378820 $Y=1061500
X2346 2359 2385 2 1 2424 2402 MUX2 $T=383160 1061880 0 0 $X=383160 $Y=1061500
X2347 2391 2398 2 1 2302 2402 MUX2 $T=383780 1041720 0 0 $X=383780 $Y=1041340
X2348 2360 2420 2 1 2285 2402 MUX2 $T=389980 1082040 0 180 $X=385640 $Y=1076620
X2349 2442 2411 2 1 2340 2402 MUX2 $T=391220 1041720 0 180 $X=386880 $Y=1036300
X2350 2414 2411 2 1 2336 2454 MUX2 $T=388120 1021560 0 0 $X=388120 $Y=1021180
X2351 2267 2465 2 1 2362 2454 MUX2 $T=397420 1031640 0 180 $X=393080 $Y=1026220
X2352 2325 2420 2 1 2216 218 MUX2 $T=393080 1071960 0 0 $X=393080 $Y=1071580
X2353 2287 2398 2 1 2346 2488 MUX2 $T=394940 1001400 0 0 $X=394940 $Y=1001020
X2354 2370 2465 2 1 2387 2402 MUX2 $T=401140 1041720 0 180 $X=396800 $Y=1036300
X2355 2369 2486 2 1 2514 2454 MUX2 $T=399900 1031640 1 0 $X=399900 $Y=1026220
X2356 2333 2465 2 1 2511 2488 MUX2 $T=399900 1041720 0 0 $X=399900 $Y=1041340
X2357 2490 2486 2 1 2443 2402 MUX2 $T=405480 1041720 0 180 $X=401140 $Y=1036300
X2358 2536 2522 2 1 2462 198 MUX2 $T=406720 1071960 1 180 $X=402380 $Y=1071580
X2359 2344 2398 2 1 2460 227 MUX2 $T=404240 1051800 1 0 $X=404240 $Y=1046380
X2360 2527 2486 2 1 2555 2488 MUX2 $T=405480 1041720 1 0 $X=405480 $Y=1036300
X2361 2521 2522 2 1 2552 2454 MUX2 $T=405480 1061880 0 0 $X=405480 $Y=1061500
X2362 2588 2522 2 1 2546 218 MUX2 $T=415400 1071960 1 180 $X=411060 $Y=1071580
X2363 2519 2465 2 1 2567 2582 MUX2 $T=418500 1041720 0 180 $X=414160 $Y=1036300
X2364 2587 2411 2 1 2608 227 MUX2 $T=414780 1051800 1 0 $X=414780 $Y=1046380
X2365 2670 240 2 1 2635 2642 MUX2 $T=427180 1071960 1 180 $X=422840 $Y=1071580
X2366 2677 2411 2 1 2629 2582 MUX2 $T=429040 1031640 1 180 $X=424700 $Y=1031260
X2367 2649 240 2 1 2685 241 MUX2 $T=424700 1061880 0 0 $X=424700 $Y=1061500
X2368 2683 2738 2 1 2623 2582 MUX2 $T=436480 1041720 0 180 $X=432140 $Y=1036300
X2369 259 205 2 1 2700 2642 MUX2 $T=438340 1082040 0 180 $X=434000 $Y=1076620
X2370 2693 260 2 1 2706 2488 MUX2 $T=439580 920760 1 180 $X=435240 $Y=920380
X2371 257 251 2 1 264 2642 MUX2 $T=435860 1082040 0 0 $X=435860 $Y=1081660
X2372 2752 2522 2 1 2699 227 MUX2 $T=443300 1071960 0 180 $X=438960 $Y=1066540
X2373 2615 2420 2 1 2755 265 MUX2 $T=439580 1071960 0 0 $X=439580 $Y=1071580
X2374 2712 266 2 1 2715 2702 MUX2 $T=445160 920760 1 180 $X=440820 $Y=920380
X2375 2713 2744 2 1 2760 267 MUX2 $T=440820 1011480 0 0 $X=440820 $Y=1011100
X2376 2745 2549 2 1 2764 2582 MUX2 $T=442060 1031640 1 0 $X=442060 $Y=1026220
X2377 272 260 2 1 2746 268 MUX2 $T=450120 920760 1 180 $X=445780 $Y=920380
X2378 2307 2645 2 1 2766 267 MUX2 $T=450120 1011480 1 180 $X=445780 $Y=1011100
X2379 269 2645 2 1 2741 2800 MUX2 $T=447020 1041720 1 0 $X=447020 $Y=1036300
X2380 2736 2738 2 1 2804 2800 MUX2 $T=447640 1051800 1 0 $X=447640 $Y=1046380
X2381 276 2385 2 1 2758 2790 MUX2 $T=452600 1071960 1 180 $X=448260 $Y=1071580
X2382 274 260 2 1 2769 267 MUX2 $T=453220 900600 1 180 $X=448880 $Y=900220
X2383 2832 2522 2 1 2788 2582 MUX2 $T=456320 1041720 0 180 $X=451980 $Y=1036300
X2384 2836 282 2 1 2791 2702 MUX2 $T=458180 920760 0 180 $X=453840 $Y=915340
X2385 2765 266 2 1 2816 268 MUX2 $T=458180 920760 1 180 $X=453840 $Y=920380
X2386 2842 2522 2 1 2821 2819 MUX2 $T=458800 1051800 0 180 $X=454460 $Y=1046380
X2387 2762 2420 2 1 2794 2819 MUX2 $T=459420 1061880 0 180 $X=455080 $Y=1056460
X2388 2873 292 2 1 2841 2642 MUX2 $T=464380 1071960 1 180 $X=460040 $Y=1071580
X2389 287 2420 2 1 2861 2582 MUX2 $T=461280 1031640 0 0 $X=461280 $Y=1031260
X2390 296 292 2 1 288 284 MUX2 $T=465620 1082040 1 180 $X=461280 $Y=1081660
X2391 2894 282 2 1 2852 270 MUX2 $T=469960 900600 1 180 $X=465620 $Y=900220
X2392 2878 282 2 1 2895 2902 MUX2 $T=465620 920760 1 0 $X=465620 $Y=915340
X2393 2905 299 2 1 2881 285 MUX2 $T=469960 1082040 1 180 $X=465620 $Y=1081660
X2394 2918 292 2 1 2897 2819 MUX2 $T=473680 1061880 0 180 $X=469340 $Y=1056460
X2395 2930 299 2 1 2909 2642 MUX2 $T=474920 1071960 1 180 $X=470580 $Y=1071580
X2396 2686 307 2 1 2964 2702 MUX2 $T=476160 920760 1 0 $X=476160 $Y=915340
X2397 2969 307 2 1 2914 2902 MUX2 $T=481120 920760 1 180 $X=476780 $Y=920380
X2398 2983 299 2 1 2953 2819 MUX2 $T=484220 1051800 1 180 $X=479880 $Y=1051420
X2399 3010 2838 2 1 2977 2992 MUX2 $T=489800 981240 0 180 $X=485460 $Y=975820
X2400 2988 2993 2 1 3015 2992 MUX2 $T=486700 1001400 1 0 $X=486700 $Y=995980
X2401 3017 3012 2 1 2934 2888 MUX2 $T=491040 1041720 0 180 $X=486700 $Y=1036300
X2402 2956 322 2 1 2998 2642 MUX2 $T=491040 1051800 1 180 $X=486700 $Y=1051420
X2403 3001 2645 2 1 3034 3023 MUX2 $T=487320 1011480 0 0 $X=487320 $Y=1011100
X2404 3028 3012 2 1 2991 285 MUX2 $T=492900 1071960 1 180 $X=488560 $Y=1071580
X2405 3006 321 2 1 3036 2902 MUX2 $T=489180 920760 0 0 $X=489180 $Y=920380
X2406 324 321 2 1 3038 2702 MUX2 $T=490420 920760 1 0 $X=490420 $Y=915340
X2407 3022 2823 2 1 3042 3023 MUX2 $T=491040 1001400 1 0 $X=491040 $Y=995980
X2408 3072 2947 2 1 3014 2992 MUX2 $T=498480 981240 0 180 $X=494140 $Y=975820
X2409 3011 2744 2 1 3061 3023 MUX2 $T=494140 1011480 0 0 $X=494140 $Y=1011100
X2410 3040 322 2 1 3065 2990 MUX2 $T=494140 1051800 1 0 $X=494140 $Y=1046380
X2411 3048 3031 2 1 3066 3067 MUX2 $T=496000 940920 0 0 $X=496000 $Y=940540
X2412 3050 2744 2 1 3068 2992 MUX2 $T=496000 951000 1 0 $X=496000 $Y=945580
X2413 3051 2823 2 1 3070 2992 MUX2 $T=496000 1001400 1 0 $X=496000 $Y=995980
X2414 2242 2948 2 1 2966 3062 MUX2 $T=499100 961080 1 0 $X=499100 $Y=955660
X2415 3064 3012 2 1 3081 2790 MUX2 $T=499100 1061880 1 0 $X=499100 $Y=1056460
X2416 3052 3012 2 1 3090 335 MUX2 $T=499720 1082040 1 0 $X=499720 $Y=1076620
X2417 338 3060 2 1 3009 331 MUX2 $T=505920 910680 0 180 $X=501580 $Y=905260
X2418 3076 3012 2 1 3092 339 MUX2 $T=501580 1071960 0 0 $X=501580 $Y=1071580
X2419 3128 3127 2 1 3098 285 MUX2 $T=510880 1071960 1 180 $X=506540 $Y=1071580
X2420 3116 3012 2 1 3135 2990 MUX2 $T=508400 1041720 0 0 $X=508400 $Y=1041340
X2421 348 3127 2 1 3147 335 MUX2 $T=510260 1071960 1 0 $X=510260 $Y=1066540
X2422 3150 3127 2 1 3103 2790 MUX2 $T=516460 1051800 1 180 $X=512120 $Y=1051420
X2423 3140 3139 2 1 3164 351 MUX2 $T=513980 910680 0 0 $X=513980 $Y=910300
X2424 3194 3190 2 1 3165 3067 MUX2 $T=523280 951000 0 180 $X=518940 $Y=945580
X2425 3187 3195 2 1 3136 335 MUX2 $T=523280 1071960 1 180 $X=518940 $Y=1071580
X2426 3215 3127 2 1 3133 2990 MUX2 $T=527620 1031640 1 180 $X=523280 $Y=1031260
X2427 3220 3195 2 1 3167 351 MUX2 $T=528860 1061880 0 180 $X=524520 $Y=1056460
X2428 2304 3169 2 1 3138 3217 MUX2 $T=525140 971160 1 0 $X=525140 $Y=965740
X2429 3225 3195 2 1 3246 2790 MUX2 $T=529480 1061880 1 0 $X=529480 $Y=1056460
X2430 3249 376 2 1 3193 3229 MUX2 $T=534440 1071960 1 180 $X=530100 $Y=1071580
X2431 3201 3195 2 1 3248 2990 MUX2 $T=530720 1041720 1 0 $X=530720 $Y=1036300
X2432 379 3127 2 1 3206 339 MUX2 $T=536300 1061880 1 180 $X=531960 $Y=1061500
X2433 3265 3127 2 1 3161 2888 MUX2 $T=537540 1041720 1 180 $X=533200 $Y=1041340
X2434 393 391 2 1 3262 3229 MUX2 $T=543120 1071960 1 180 $X=538780 $Y=1071580
X2435 3298 401 2 1 3278 2902 MUX2 $T=548080 920760 0 180 $X=543740 $Y=915340
X2436 3292 3195 2 1 3338 3276 MUX2 $T=544980 1051800 1 0 $X=544980 $Y=1046380
X2437 405 401 2 1 398 294 MUX2 $T=549940 900600 1 180 $X=545600 $Y=900220
X2438 3352 3354 2 1 3312 402 MUX2 $T=552420 1071960 0 180 $X=548080 $Y=1066540
X2439 3337 3321 2 1 3261 3217 MUX2 $T=553660 981240 0 180 $X=549320 $Y=975820
X2440 2339 3353 2 1 3279 3217 MUX2 $T=553660 991320 1 180 $X=549320 $Y=990940
X2441 414 3358 2 1 417 294 MUX2 $T=553040 900600 0 0 $X=553040 $Y=900220
X2442 418 3373 2 1 3286 3359 MUX2 $T=557380 961080 0 180 $X=553040 $Y=955660
X2443 3351 3369 2 1 3403 3217 MUX2 $T=556140 991320 0 0 $X=556140 $Y=990940
X2444 3375 3354 2 1 3360 339 MUX2 $T=561100 1061880 1 180 $X=556760 $Y=1061500
X2445 3349 412 2 1 3313 3229 MUX2 $T=561100 1082040 0 180 $X=556760 $Y=1076620
X2446 3363 3290 2 1 3389 3067 MUX2 $T=557380 940920 0 0 $X=557380 $Y=940540
X2447 420 3358 2 1 3419 383 MUX2 $T=558000 910680 1 0 $X=558000 $Y=905260
X2448 3411 3417 2 1 3346 392 MUX2 $T=562340 1051800 1 180 $X=558000 $Y=1051420
X2449 430 431 2 1 424 402 MUX2 $T=564820 1082040 1 180 $X=560480 $Y=1081660
X2450 3402 3358 2 1 3421 3053 MUX2 $T=561100 920760 1 0 $X=561100 $Y=915340
X2451 3405 3414 2 1 3431 3067 MUX2 $T=561720 940920 0 0 $X=561720 $Y=940540
X2452 3451 401 2 1 3427 3053 MUX2 $T=569780 920760 0 180 $X=565440 $Y=915340
X2453 441 3417 2 1 3444 339 MUX2 $T=572260 1071960 1 180 $X=567920 $Y=1071580
X2454 3474 431 2 1 3446 3229 MUX2 $T=574120 1082040 0 180 $X=569780 $Y=1076620
X2455 3438 3354 2 1 3491 3276 MUX2 $T=572260 1051800 0 0 $X=572260 $Y=1051420
X2456 449 3353 2 1 3450 3023 MUX2 $T=577220 1021560 1 180 $X=572880 $Y=1021180
X2457 3467 3417 2 1 3488 402 MUX2 $T=572880 1061880 0 0 $X=572880 $Y=1061500
X2458 3485 455 2 1 3489 3053 MUX2 $T=581560 920760 0 180 $X=577220 $Y=915340
X2459 462 3354 2 1 3475 2790 MUX2 $T=581560 1061880 1 180 $X=577220 $Y=1061500
X2460 3508 455 2 1 3479 3401 MUX2 $T=582800 930840 0 180 $X=578460 $Y=925420
X2461 458 3354 2 1 3502 3229 MUX2 $T=580940 1051800 0 0 $X=580940 $Y=1051420
X2462 3543 3417 2 1 456 460 MUX2 $T=585900 1082040 1 180 $X=581560 $Y=1081660
X2463 466 455 2 1 472 383 MUX2 $T=582800 900600 0 0 $X=582800 $Y=900220
X2464 468 3354 2 1 3547 3548 MUX2 $T=584660 1061880 0 0 $X=584660 $Y=1061500
X2465 3533 3378 2 1 3549 3023 MUX2 $T=585900 1021560 1 0 $X=585900 $Y=1016140
X2466 3540 3417 2 1 3551 3229 MUX2 $T=586520 1051800 0 0 $X=586520 $Y=1051420
X2467 3241 3290 2 1 3576 483 MUX2 $T=592720 940920 0 0 $X=592720 $Y=940540
X2468 3561 482 2 1 3580 3492 MUX2 $T=593340 920760 1 0 $X=593340 $Y=915340
X2469 3538 3290 2 1 3566 3587 MUX2 $T=595200 1011480 0 0 $X=595200 $Y=1011100
X2470 493 3586 2 1 3578 485 MUX2 $T=602020 951000 0 180 $X=597680 $Y=945580
X2471 490 3586 2 1 3605 483 MUX2 $T=600780 961080 1 0 $X=600780 $Y=955660
X2472 2524 3290 2 1 3622 3629 MUX2 $T=600780 971160 1 0 $X=600780 $Y=965740
X2473 492 3290 2 1 3617 485 MUX2 $T=601400 940920 0 0 $X=601400 $Y=940540
X2474 488 3378 2 1 3632 3629 MUX2 $T=602020 981240 0 0 $X=602020 $Y=980860
X2475 3630 498 2 1 3560 494 MUX2 $T=606980 1082040 1 180 $X=602640 $Y=1081660
X2476 503 482 2 1 3601 3401 MUX2 $T=609460 920760 1 180 $X=605120 $Y=920380
X2477 3591 3644 2 1 3553 3616 MUX2 $T=610080 1061880 0 180 $X=605740 $Y=1056460
X2478 3648 3647 2 1 3567 3401 MUX2 $T=610700 1041720 0 180 $X=606360 $Y=1036300
X2479 506 498 2 1 500 501 MUX2 $T=611320 1082040 1 180 $X=606980 $Y=1081660
X2480 3651 504 2 1 3626 3492 MUX2 $T=611940 910680 0 180 $X=607600 $Y=905260
X2481 3624 502 2 1 3653 3548 MUX2 $T=607600 1082040 1 0 $X=607600 $Y=1076620
X2482 512 3657 2 1 3579 3359 MUX2 $T=613180 971160 0 180 $X=608840 $Y=965740
X2483 3645 504 2 1 3662 3556 MUX2 $T=609460 920760 0 0 $X=609460 $Y=920380
X2484 3608 3677 2 1 3604 3616 MUX2 $T=615660 1021560 1 180 $X=611320 $Y=1021180
X2485 3680 3684 2 1 3593 3616 MUX2 $T=616280 1041720 0 180 $X=611940 $Y=1036300
X2486 3683 3682 2 1 3658 3616 MUX2 $T=616280 1061880 0 180 $X=611940 $Y=1056460
X2487 3686 3679 2 1 3581 3654 MUX2 $T=616900 991320 1 180 $X=612560 $Y=990940
X2488 519 3647 2 1 3597 3654 MUX2 $T=617520 1001400 1 180 $X=613180 $Y=1001020
X2489 513 3647 2 1 3585 3687 MUX2 $T=613180 1031640 1 0 $X=613180 $Y=1026220
X2490 3661 3644 2 1 3575 3697 MUX2 $T=613180 1041720 0 0 $X=613180 $Y=1041340
X2491 3665 504 2 1 3698 3401 MUX2 $T=613800 920760 0 0 $X=613800 $Y=920380
X2492 3649 518 2 1 3668 517 MUX2 $T=618760 910680 0 180 $X=614420 $Y=905260
X2493 2625 518 2 1 3716 3556 MUX2 $T=616900 920760 1 0 $X=616900 $Y=915340
X2494 3719 3702 2 1 3655 3359 MUX2 $T=621860 971160 0 180 $X=617520 $Y=965740
X2495 3695 3684 2 1 3720 3687 MUX2 $T=617520 1021560 0 0 $X=617520 $Y=1021180
X2496 3740 3726 2 1 3667 3708 MUX2 $T=623100 940920 1 180 $X=618760 $Y=940540
X2497 3712 502 2 1 3732 501 MUX2 $T=619380 1082040 1 0 $X=619380 $Y=1076620
X2498 3742 3684 2 1 3717 3697 MUX2 $T=624960 1041720 0 180 $X=620620 $Y=1036300
X2499 3568 3704 2 1 3749 3654 MUX2 $T=621240 1011480 1 0 $X=621240 $Y=1006060
X2500 528 518 2 1 3772 3722 MUX2 $T=621860 920760 1 0 $X=621860 $Y=915340
X2501 3750 3752 2 1 3631 3708 MUX2 $T=626200 951000 0 180 $X=621860 $Y=945580
X2502 3640 3677 2 1 3763 3620 MUX2 $T=624340 1031640 0 0 $X=624340 $Y=1031260
X2503 3767 3644 2 1 3707 3747 MUX2 $T=629300 1061880 1 180 $X=624960 $Y=1061500
X2504 3780 3752 2 1 3755 485 MUX2 $T=631160 940920 1 180 $X=626820 $Y=940540
X2505 538 3677 2 1 3705 3747 MUX2 $T=631780 1021560 0 180 $X=627440 $Y=1016140
X2506 3770 3644 2 1 3779 543 MUX2 $T=629300 1061880 0 0 $X=629300 $Y=1061500
X2507 3782 3677 2 1 3804 3697 MUX2 $T=632400 1041720 1 0 $X=632400 $Y=1036300
X2508 551 544 2 1 541 3722 MUX2 $T=638600 910680 0 180 $X=634260 $Y=905260
X2509 3797 544 2 1 3811 3556 MUX2 $T=636120 920760 0 0 $X=636120 $Y=920380
X2510 558 3684 2 1 3805 3747 MUX2 $T=642320 1031640 0 180 $X=637980 $Y=1026220
X2511 3823 3682 2 1 3807 543 MUX2 $T=642320 1061880 0 180 $X=637980 $Y=1056460
X2512 3845 544 2 1 3798 557 MUX2 $T=646040 920760 1 180 $X=641700 $Y=920380
X2513 3833 3657 2 1 3775 3852 MUX2 $T=643560 1082040 1 0 $X=643560 $Y=1076620
X2514 3847 3677 2 1 3862 3806 MUX2 $T=646660 1041720 1 0 $X=646660 $Y=1036300
X2515 3864 568 2 1 3809 557 MUX2 $T=651620 920760 1 180 $X=647280 $Y=920380
X2516 3663 546 2 1 3885 483 MUX2 $T=647900 940920 0 0 $X=647900 $Y=940540
X2517 3614 3677 2 1 3835 3863 MUX2 $T=647900 1031640 0 0 $X=647900 $Y=1031260
X2518 3871 3702 2 1 3837 3852 MUX2 $T=652240 1082040 0 180 $X=647900 $Y=1076620
X2519 3889 3644 2 1 3849 3863 MUX2 $T=654720 1061880 0 180 $X=650380 $Y=1056460
X2520 3887 3795 2 1 3817 3629 MUX2 $T=655340 961080 0 180 $X=651000 $Y=955660
X2521 575 568 2 1 3909 3854 MUX2 $T=652860 920760 1 0 $X=652860 $Y=915340
X2522 3893 568 2 1 3924 3722 MUX2 $T=655960 910680 1 0 $X=655960 $Y=905260
X2523 3762 3839 2 1 3861 3629 MUX2 $T=661540 981240 1 180 $X=657200 $Y=980860
X2524 591 546 2 1 3905 3629 MUX2 $T=662160 961080 0 180 $X=657820 $Y=955660
X2525 3915 3684 2 1 3935 3863 MUX2 $T=659060 1031640 0 0 $X=659060 $Y=1031260
X2526 3920 546 2 1 3939 3852 MUX2 $T=659680 1071960 0 0 $X=659680 $Y=1071580
X2527 3956 3858 2 1 3986 3987 MUX2 $T=665880 1031640 0 0 $X=665880 $Y=1031260
X2528 3973 3860 2 1 4002 3969 MUX2 $T=668360 1041720 0 0 $X=668360 $Y=1041340
X2529 3943 3839 2 1 4004 3987 MUX2 $T=668980 1021560 1 0 $X=668980 $Y=1016140
X2530 609 606 2 1 603 3852 MUX2 $T=673320 1082040 1 180 $X=668980 $Y=1081660
X2531 604 3812 2 1 4006 3852 MUX2 $T=669600 1082040 1 0 $X=669600 $Y=1076620
X2532 4016 616 2 1 3974 557 MUX2 $T=675800 920760 1 180 $X=671460 $Y=920380
X2533 3637 605 2 1 3950 607 MUX2 $T=677040 940920 1 180 $X=672700 $Y=940540
X2534 622 605 2 1 613 3852 MUX2 $T=678900 1082040 1 180 $X=674560 $Y=1081660
X2535 3979 616 2 1 3929 3854 MUX2 $T=679520 920760 0 180 $X=675180 $Y=915340
X2536 3988 3975 2 1 4027 620 MUX2 $T=681380 940920 1 180 $X=677040 $Y=940540
X2537 623 616 2 1 3957 3722 MUX2 $T=678900 910680 1 0 $X=678900 $Y=905260
X2538 631 4061 2 1 3953 3987 MUX2 $T=683240 1051800 1 180 $X=678900 $Y=1051420
X2539 4045 4055 2 1 4056 4033 MUX2 $T=682620 991320 1 0 $X=682620 $Y=985900
X2540 636 4055 2 1 4022 3587 MUX2 $T=686960 1011480 1 180 $X=682620 $Y=1011100
X2541 4096 4088 2 1 4068 4033 MUX2 $T=688200 971160 0 180 $X=683860 $Y=965740
X2542 642 4086 2 1 4035 3987 MUX2 $T=688200 1051800 1 180 $X=683860 $Y=1051420
X2543 4090 4088 2 1 4026 3969 MUX2 $T=688200 1071960 1 180 $X=683860 $Y=1071580
X2544 4007 634 2 1 4106 3854 MUX2 $T=684480 920760 0 0 $X=684480 $Y=920380
X2545 4077 4066 2 1 4105 4033 MUX2 $T=684480 1001400 1 0 $X=684480 $Y=995980
X2546 4073 4066 2 1 4097 3987 MUX2 $T=684480 1031640 0 0 $X=684480 $Y=1031260
X2547 4111 4055 2 1 4042 4054 MUX2 $T=691300 991320 0 180 $X=686960 $Y=985900
X2548 4017 4087 2 1 4119 4054 MUX2 $T=687580 961080 1 0 $X=687580 $Y=955660
X2549 4122 4086 2 1 4099 3620 MUX2 $T=692540 1051800 1 180 $X=688200 $Y=1051420
X2550 4104 4086 2 1 4110 4033 MUX2 $T=689440 1011480 0 0 $X=689440 $Y=1011100
X2551 4112 648 2 1 645 567 MUX2 $T=695640 1082040 1 180 $X=691300 $Y=1081660
X2552 4118 4066 2 1 4144 3620 MUX2 $T=691920 1031640 1 0 $X=691920 $Y=1026220
X2553 4013 4061 2 1 4121 3620 MUX2 $T=696880 1051800 1 180 $X=692540 $Y=1051420
X2554 3985 4141 2 1 4102 4033 MUX2 $T=697500 1011480 0 180 $X=693160 $Y=1006060
X2555 4037 4149 2 1 4129 3620 MUX2 $T=697500 1041720 0 180 $X=693160 $Y=1036300
X2556 4155 4151 2 1 4107 4131 MUX2 $T=698740 1071960 1 180 $X=694400 $Y=1071580
X2557 647 4087 2 1 4152 4033 MUX2 $T=695020 971160 0 0 $X=695020 $Y=970780
X2558 4135 634 2 1 4169 4180 MUX2 $T=698120 920760 0 0 $X=698120 $Y=920380
X2559 4202 660 2 1 4182 4114 MUX2 $T=706800 920760 0 180 $X=702460 $Y=915340
X2560 4206 4149 2 1 4163 4103 MUX2 $T=706800 1031640 1 180 $X=702460 $Y=1031260
X2561 4179 661 2 1 4187 4132 MUX2 $T=707420 910680 0 180 $X=703080 $Y=905260
X2562 4209 4086 2 1 4189 4103 MUX2 $T=707420 1051800 1 180 $X=703080 $Y=1051420
X2563 3933 661 2 1 4160 4114 MUX2 $T=708040 920760 1 180 $X=703700 $Y=920380
X2564 4215 655 2 1 654 567 MUX2 $T=708040 1082040 0 180 $X=703700 $Y=1076620
X2565 4084 4061 2 1 4186 4103 MUX2 $T=709900 1061880 1 180 $X=705560 $Y=1061500
X2566 4229 4230 2 1 4201 4103 MUX2 $T=711140 1031640 1 180 $X=706800 $Y=1031260
X2567 4218 4149 2 1 4210 3747 MUX2 $T=713620 1021560 0 180 $X=709280 $Y=1016140
X2568 4136 661 2 1 4257 4180 MUX2 $T=711760 920760 0 0 $X=711760 $Y=920380
X2569 4245 3975 2 1 4258 483 MUX2 $T=713620 940920 0 0 $X=713620 $Y=940540
X2570 4220 4230 2 1 4196 3806 MUX2 $T=718580 1031640 1 180 $X=714240 $Y=1031260
X2571 677 4061 2 1 4239 667 MUX2 $T=720440 1041720 1 180 $X=716100 $Y=1041340
X2572 4280 4086 2 1 4244 667 MUX2 $T=721060 1061880 0 180 $X=716720 $Y=1056460
X2573 671 4230 2 1 4283 667 MUX2 $T=717960 1011480 0 0 $X=717960 $Y=1011100
X2574 4261 648 2 1 682 680 MUX2 $T=717960 1082040 0 0 $X=717960 $Y=1081660
X2575 4262 660 2 1 4293 4180 MUX2 $T=718580 920760 1 0 $X=718580 $Y=915340
X2576 674 660 2 1 4294 4132 MUX2 $T=719820 910680 1 0 $X=719820 $Y=905260
X2577 4251 655 2 1 4317 680 MUX2 $T=719820 1082040 1 0 $X=719820 $Y=1076620
X2578 4314 4308 2 1 4276 3806 MUX2 $T=726020 1041720 0 180 $X=721680 $Y=1036300
X2579 4347 4357 2 1 4319 3806 MUX2 $T=730980 1041720 0 180 $X=726640 $Y=1036300
X2580 4351 696 2 1 4383 4114 MUX2 $T=732220 920760 1 0 $X=732220 $Y=915340
X2581 4358 696 2 1 4373 4180 MUX2 $T=732220 930840 1 0 $X=732220 $Y=925420
X2582 698 4230 2 1 4388 4378 MUX2 $T=733460 1021560 0 0 $X=733460 $Y=1021180
X2583 4371 644 2 1 4390 680 MUX2 $T=734080 1082040 0 0 $X=734080 $Y=1081660
X2584 4391 4230 2 1 4409 4413 MUX2 $T=737800 1021560 0 0 $X=737800 $Y=1021180
X2585 4392 706 2 1 4417 4180 MUX2 $T=738420 920760 0 0 $X=738420 $Y=920380
X2586 4396 706 2 1 4414 4132 MUX2 $T=739040 910680 0 0 $X=739040 $Y=910300
X2587 4397 701 2 1 4416 709 MUX2 $T=739040 1082040 0 0 $X=739040 $Y=1081660
X2588 712 706 2 1 4395 705 MUX2 $T=744620 900600 1 180 $X=740280 $Y=900220
X2589 4404 706 2 1 4420 4114 MUX2 $T=740900 920760 1 0 $X=740900 $Y=915340
X2590 708 4149 2 1 4428 4413 MUX2 $T=742760 1031640 0 0 $X=742760 $Y=1031260
X2591 713 696 2 1 4433 4132 MUX2 $T=744620 920760 0 0 $X=744620 $Y=920380
X2592 4419 4357 2 1 4435 4413 MUX2 $T=744620 1061880 0 0 $X=744620 $Y=1061500
X2593 4437 4357 2 1 4440 711 MUX2 $T=748960 1051800 0 0 $X=748960 $Y=1051420
X2594 4462 4461 2 1 4429 4441 MUX2 $T=753920 961080 0 180 $X=749580 $Y=955660
X2595 725 4446 2 1 4412 4413 MUX2 $T=755780 1021560 0 180 $X=751440 $Y=1016140
X2596 4477 4461 2 1 4436 4378 MUX2 $T=756400 981240 0 180 $X=752060 $Y=975820
X2597 4445 4461 2 1 4426 723 MUX2 $T=757020 940920 1 180 $X=752680 $Y=940540
X2598 4481 4446 2 1 4427 4454 MUX2 $T=757640 991320 1 180 $X=753300 $Y=990940
X2599 728 727 2 1 4474 709 MUX2 $T=759500 1082040 0 180 $X=755160 $Y=1076620
X2600 4507 727 2 1 4471 711 MUX2 $T=761980 1071960 0 180 $X=757640 $Y=1066540
X2601 729 4505 2 1 4465 4378 MUX2 $T=762600 981240 0 180 $X=758260 $Y=975820
X2602 4447 4505 2 1 4457 4432 MUX2 $T=762600 991320 1 180 $X=758260 $Y=990940
X2603 4519 732 2 1 4488 709 MUX2 $T=763840 1082040 0 180 $X=759500 $Y=1076620
X2604 4039 4446 2 1 4499 4132 MUX2 $T=765080 991320 0 180 $X=760740 $Y=985900
X2605 4496 735 2 1 4479 4180 MUX2 $T=765700 910680 0 180 $X=761360 $Y=905260
X2606 741 4505 2 1 4515 4454 MUX2 $T=766940 991320 1 180 $X=762600 $Y=990940
X2607 4535 4513 2 1 4443 4131 MUX2 $T=766940 1061880 0 180 $X=762600 $Y=1056460
X2608 736 4513 2 1 4467 4542 MUX2 $T=765080 1051800 0 0 $X=765080 $Y=1051420
X2609 4464 4446 2 1 4469 4545 MUX2 $T=766320 961080 0 0 $X=766320 $Y=960700
X2610 742 732 2 1 4563 711 MUX2 $T=766940 1071960 0 0 $X=766940 $Y=1071580
X2611 743 4522 2 1 4570 4131 MUX2 $T=767560 1061880 0 0 $X=767560 $Y=1061500
X2612 4556 4522 2 1 4589 4542 MUX2 $T=770040 1051800 0 0 $X=770040 $Y=1051420
X2613 4521 4539 2 1 4626 4545 MUX2 $T=776860 961080 1 0 $X=776860 $Y=955660
X2614 761 4505 2 1 4527 4623 MUX2 $T=776860 991320 0 0 $X=776860 $Y=990940
X2615 4640 781 2 1 4595 4545 MUX2 $T=783680 910680 1 180 $X=779340 $Y=910300
X2616 765 4518 2 1 4662 775 MUX2 $T=780580 930840 1 0 $X=780580 $Y=925420
X2617 771 4547 2 1 4645 775 MUX2 $T=781820 940920 1 0 $X=781820 $Y=935500
X2618 4619 4637 2 1 4660 4623 MUX2 $T=781820 991320 0 0 $X=781820 $Y=990940
X2619 4641 4637 2 1 4674 4432 MUX2 $T=783060 1001400 0 0 $X=783060 $Y=1001020
X2620 4667 4637 2 1 4642 4413 MUX2 $T=787400 1011480 1 180 $X=783060 $Y=1011100
X2621 4655 4637 2 1 4629 4545 MUX2 $T=788020 971160 0 180 $X=783680 $Y=965740
X2622 4659 4637 2 1 4683 4454 MUX2 $T=785540 981240 0 0 $X=785540 $Y=980860
X2623 4651 788 2 1 4669 4673 MUX2 $T=791740 1071960 0 180 $X=787400 $Y=1066540
X2624 792 788 2 1 4670 782 MUX2 $T=791740 1082040 0 180 $X=787400 $Y=1076620
X2625 4658 803 2 1 4666 4545 MUX2 $T=795460 920760 0 180 $X=791120 $Y=915340
X2626 4731 4709 2 1 4646 4131 MUX2 $T=796080 1071960 0 180 $X=791740 $Y=1066540
X2627 4665 4637 2 1 4671 4533 MUX2 $T=797320 961080 1 180 $X=792980 $Y=960700
X2628 809 805 2 1 4722 4717 MUX2 $T=798560 910680 0 180 $X=794220 $Y=905260
X2629 4583 4729 2 1 4754 4703 MUX2 $T=794840 971160 1 0 $X=794840 $Y=965740
X2630 806 805 2 1 4767 4761 MUX2 $T=796080 920760 1 0 $X=796080 $Y=915340
X2631 4745 4695 2 1 4712 4609 MUX2 $T=802900 971160 1 180 $X=798560 $Y=970780
X2632 817 818 2 1 4759 4673 MUX2 $T=804140 1082040 0 180 $X=799800 $Y=1076620
X2633 4534 4795 2 1 4725 4454 MUX2 $T=805380 991320 0 180 $X=801040 $Y=985900
X2634 4801 4709 2 1 4768 4542 MUX2 $T=806000 1061880 0 180 $X=801660 $Y=1056460
X2635 4538 4729 2 1 4807 4533 MUX2 $T=802900 961080 1 0 $X=802900 $Y=955660
X2636 4785 803 2 1 4810 4761 MUX2 $T=803520 910680 0 0 $X=803520 $Y=910300
X2637 4814 4795 2 1 4764 4432 MUX2 $T=807860 1001400 1 180 $X=803520 $Y=1001020
X2638 4796 4795 2 1 4836 4623 MUX2 $T=805380 991320 1 0 $X=805380 $Y=985900
X2639 4833 821 2 1 4773 4673 MUX2 $T=809720 1082040 0 180 $X=805380 $Y=1076620
X2640 4819 4795 2 1 4862 782 MUX2 $T=808480 1001400 0 0 $X=808480 $Y=1001020
X2641 4834 803 2 1 4846 829 MUX2 $T=809720 910680 1 0 $X=809720 $Y=905260
X2642 4840 4795 2 1 4857 4609 MUX2 $T=810340 991320 1 0 $X=810340 $Y=985900
X2643 4849 4695 2 1 4876 4635 MUX2 $T=812200 971160 0 0 $X=812200 $Y=970780
X2644 4855 4803 2 1 4882 4635 MUX2 $T=813440 971160 1 0 $X=813440 $Y=965740
X2645 4864 4853 2 1 4891 4761 MUX2 $T=814680 1011480 1 0 $X=814680 $Y=1006060
X2646 4892 4884 2 1 4867 4542 MUX2 $T=819020 1051800 1 180 $X=814680 $Y=1051420
X2647 4895 821 2 1 4917 850 MUX2 $T=819640 1082040 1 0 $X=819640 $Y=1076620
X2648 4906 847 2 1 4925 782 MUX2 $T=822120 910680 1 0 $X=822120 $Y=905260
X2649 4930 851 2 1 4913 829 MUX2 $T=827700 920760 0 180 $X=823360 $Y=915340
X2650 4932 4872 2 1 4899 4761 MUX2 $T=827700 1011480 1 180 $X=823360 $Y=1011100
X2651 4945 4923 2 1 4921 4911 MUX2 $T=830800 1051800 1 180 $X=826460 $Y=1051420
X2652 4949 4952 2 1 4898 4609 MUX2 $T=832040 981240 1 180 $X=827700 $Y=980860
X2653 4956 4952 2 1 4936 4432 MUX2 $T=833280 1001400 0 180 $X=828940 $Y=995980
X2654 855 4884 2 1 4958 4934 MUX2 $T=828940 1061880 1 0 $X=828940 $Y=1056460
X2655 4980 4961 2 1 4928 4955 MUX2 $T=837000 961080 1 180 $X=832660 $Y=960700
X2656 4681 4961 2 1 4979 4609 MUX2 $T=833280 951000 1 0 $X=833280 $Y=945580
X2657 4981 4952 2 1 4948 4623 MUX2 $T=837620 1001400 0 180 $X=833280 $Y=995980
X2658 4989 805 2 1 4939 4114 MUX2 $T=838240 910680 1 180 $X=833900 $Y=910300
X2659 4777 4967 2 1 4943 4955 MUX2 $T=840100 951000 1 180 $X=835760 $Y=950620
X2660 4973 4977 2 1 4991 4761 MUX2 $T=835760 1021560 0 0 $X=835760 $Y=1021180
X2661 4999 5000 2 1 4912 4432 MUX2 $T=841340 991320 1 180 $X=837000 $Y=990940
X2662 866 4933 2 1 4996 4955 MUX2 $T=838860 910680 1 0 $X=838860 $Y=905260
X2663 5017 5000 2 1 4988 4609 MUX2 $T=843200 981240 1 180 $X=838860 $Y=980860
X2664 867 864 2 1 5013 871 MUX2 $T=838860 1082040 1 0 $X=838860 $Y=1076620
X2665 5023 4977 2 1 4985 4911 MUX2 $T=844440 1041720 1 180 $X=840100 $Y=1041340
X2666 870 864 2 1 4929 868 MUX2 $T=844440 1082040 1 180 $X=840100 $Y=1081660
X2667 4812 4967 2 1 5016 5034 MUX2 $T=841340 961080 0 0 $X=841340 $Y=960700
X2668 5035 4977 2 1 4975 4934 MUX2 $T=846920 1071960 0 180 $X=842580 $Y=1066540
X2669 877 4933 2 1 5019 5018 MUX2 $T=848160 930840 0 180 $X=843820 $Y=925420
X2670 5044 5032 2 1 5022 4761 MUX2 $T=848160 1011480 1 180 $X=843820 $Y=1011100
X2671 5056 4961 2 1 5011 5034 MUX2 $T=850640 961080 1 180 $X=846300 $Y=960700
X2672 881 880 2 1 876 850 MUX2 $T=851260 1082040 1 180 $X=846920 $Y=1081660
X2673 5043 4967 2 1 5073 5018 MUX2 $T=847540 940920 0 0 $X=847540 $Y=940540
X2674 5053 5000 2 1 5075 5081 MUX2 $T=849400 981240 0 0 $X=849400 $Y=980860
X2675 5080 5095 2 1 5061 4911 MUX2 $T=854980 1041720 0 180 $X=850640 $Y=1036300
X2676 5087 5000 2 1 5033 829 MUX2 $T=855600 991320 0 180 $X=851260 $Y=985900
X2677 5092 851 2 1 5024 5070 MUX2 $T=856840 920760 0 180 $X=852500 $Y=915340
X2678 5071 5000 2 1 5040 4454 MUX2 $T=857460 1001400 0 180 $X=853120 $Y=995980
X2679 5084 851 2 1 5025 894 MUX2 $T=854980 910680 1 0 $X=854980 $Y=905260
X2680 895 851 2 1 5060 5086 MUX2 $T=859320 920760 1 180 $X=854980 $Y=920380
X2681 5102 5095 2 1 5106 4934 MUX2 $T=856840 1061880 0 0 $X=856840 $Y=1061500
X2682 889 880 2 1 5097 871 MUX2 $T=856840 1071960 0 0 $X=856840 $Y=1071580
X2683 5122 5114 2 1 5105 829 MUX2 $T=861800 991320 0 180 $X=857460 $Y=985900
X2684 5127 5138 2 1 5093 829 MUX2 $T=862420 951000 1 180 $X=858080 $Y=950620
X2685 5121 5109 2 1 5103 829 MUX2 $T=862420 971160 1 180 $X=858080 $Y=970780
X2686 4986 4933 2 1 5145 5086 MUX2 $T=859940 920760 0 0 $X=859940 $Y=920380
X2687 5113 5108 2 1 5151 5070 MUX2 $T=859940 940920 0 0 $X=859940 $Y=940540
X2688 5133 5138 2 1 5038 5070 MUX2 $T=864280 951000 0 180 $X=859940 $Y=945580
X2689 5150 5114 2 1 5117 5070 MUX2 $T=866140 1001400 0 180 $X=861800 $Y=995980
X2690 898 4933 2 1 5160 894 MUX2 $T=863660 910680 1 0 $X=863660 $Y=905260
X2691 908 5109 2 1 5152 4703 MUX2 $T=871720 961080 1 180 $X=867380 $Y=960700
X2692 5194 909 2 1 5139 871 MUX2 $T=871720 1071960 0 180 $X=867380 $Y=1066540
X2693 5170 5149 2 1 5189 4934 MUX2 $T=868620 1061880 0 0 $X=868620 $Y=1061500
X2694 5211 5114 2 1 5157 5176 MUX2 $T=874200 981240 1 180 $X=869860 $Y=980860
X2695 5208 911 2 1 5153 5086 MUX2 $T=875440 920760 0 180 $X=871100 $Y=915340
X2696 5201 4967 2 1 5163 4635 MUX2 $T=875440 951000 0 180 $X=871100 $Y=945580
X2697 5229 911 2 1 5178 4955 MUX2 $T=879160 910680 1 180 $X=874820 $Y=910300
X2698 5217 5108 2 1 5241 4635 MUX2 $T=876060 951000 1 0 $X=876060 $Y=945580
X2699 5238 917 2 1 5218 871 MUX2 $T=880400 1071960 0 180 $X=876060 $Y=1066540
X2700 5219 909 2 1 5207 868 MUX2 $T=876060 1082040 0 0 $X=876060 $Y=1081660
X2701 5197 5224 2 1 5247 5176 MUX2 $T=877300 981240 0 0 $X=877300 $Y=980860
X2702 5232 5109 2 1 5282 5258 MUX2 $T=879160 971160 1 0 $X=879160 $Y=965740
X2703 5237 911 2 1 5261 5018 MUX2 $T=879780 920760 0 0 $X=879780 $Y=920380
X2704 5273 5138 2 1 5246 4533 MUX2 $T=885360 951000 1 180 $X=881020 $Y=950620
X2705 5260 5263 2 1 5272 5262 MUX2 $T=882880 991320 0 0 $X=882880 $Y=990940
X2706 5289 5300 2 1 5216 4934 MUX2 $T=887840 1061880 1 180 $X=883500 $Y=1061500
X2707 5317 5284 2 1 5283 5262 MUX2 $T=891560 1001400 0 180 $X=887220 $Y=995980
X2708 5314 5245 2 1 5335 4911 MUX2 $T=890320 1061880 0 0 $X=890320 $Y=1061500
X2709 5337 847 2 1 5308 5086 MUX2 $T=895280 920760 0 180 $X=890940 $Y=915340
X2710 5326 847 2 1 5344 4955 MUX2 $T=892800 910680 0 0 $X=892800 $Y=910300
X2711 5349 5149 2 1 5310 4911 MUX2 $T=897140 1051800 1 180 $X=892800 $Y=1051420
X2712 5339 847 2 1 5362 5018 MUX2 $T=895280 920760 1 0 $X=895280 $Y=915340
X2713 5348 5300 2 1 5387 4911 MUX2 $T=899000 1051800 1 0 $X=899000 $Y=1046380
X2714 5389 5372 2 1 5364 5258 MUX2 $T=903960 971160 1 180 $X=899620 $Y=970780
X2715 5388 956 2 1 5373 5018 MUX2 $T=905820 920760 0 180 $X=901480 $Y=915340
X2716 954 941 2 1 5366 5395 MUX2 $T=902720 1071960 0 0 $X=902720 $Y=1071580
X2717 5329 956 2 1 5405 4955 MUX2 $T=904580 910680 1 0 $X=904580 $Y=905260
X2718 961 956 2 1 5414 906 MUX2 $T=905820 900600 0 0 $X=905820 $Y=900220
X2719 5390 956 2 1 5418 948 MUX2 $T=905820 920760 1 0 $X=905820 $Y=915340
X2720 962 941 2 1 967 868 MUX2 $T=906440 1082040 1 0 $X=906440 $Y=1076620
X2721 5445 5442 2 1 5381 5433 MUX2 $T=919460 1051800 1 180 $X=915120 $Y=1051420
X2722 5448 5442 2 1 5382 971 MUX2 $T=921320 1061880 1 180 $X=916980 $Y=1061500
X2723 5434 972 2 1 5455 5433 MUX2 $T=916980 1082040 1 0 $X=916980 $Y=1076620
X2724 5441 5415 2 1 5464 5258 MUX2 $T=918220 981240 0 0 $X=918220 $Y=980860
X2725 5470 5457 2 1 5409 485 MUX2 $T=923180 940920 0 180 $X=918840 $Y=935500
X2726 980 5452 2 1 5469 970 MUX2 $T=920700 1041720 1 0 $X=920700 $Y=1036300
X2727 995 5452 2 1 5404 5395 MUX2 $T=926900 1041720 1 180 $X=922560 $Y=1041340
X2728 997 999 2 1 5479 987 MUX2 $T=928140 920760 1 180 $X=923800 $Y=920380
X2729 5428 5452 2 1 5481 5433 MUX2 $T=928140 1061880 0 180 $X=923800 $Y=1056460
X2730 5480 5442 2 1 5489 5262 MUX2 $T=928760 1031640 1 180 $X=924420 $Y=1031260
X2731 5492 991 2 1 5509 5433 MUX2 $T=925660 1082040 0 0 $X=925660 $Y=1081660
X2732 5518 5490 2 1 5473 5498 MUX2 $T=930620 940920 0 180 $X=926280 $Y=935500
X2733 5513 5457 2 1 5468 5496 MUX2 $T=931240 951000 0 180 $X=926900 $Y=945580
X2734 1002 5508 2 1 5419 5500 MUX2 $T=931860 1011480 0 180 $X=927520 $Y=1006060
X2735 5540 5508 2 1 5440 5176 MUX2 $T=933720 1011480 1 180 $X=929380 $Y=1011100
X2736 1004 5523 2 1 5549 5500 MUX2 $T=931860 1011480 1 0 $X=931860 $Y=1006060
X2737 5516 5537 2 1 5524 987 MUX2 $T=936820 920760 1 180 $X=932480 $Y=920380
X2738 5554 5527 2 1 5510 5496 MUX2 $T=937440 961080 1 180 $X=933100 $Y=960700
X2739 5555 5523 2 1 5449 5176 MUX2 $T=937440 1021560 0 180 $X=933100 $Y=1016140
X2740 5511 5452 2 1 5551 5262 MUX2 $T=933720 1031640 0 0 $X=933720 $Y=1031260
X2741 5542 5537 2 1 5568 5496 MUX2 $T=934960 951000 0 0 $X=934960 $Y=950620
X2742 5580 1018 2 1 5478 987 MUX2 $T=941160 910680 0 180 $X=936820 $Y=905260
X2743 5506 5537 2 1 5581 5576 MUX2 $T=936820 930840 1 0 $X=936820 $Y=925420
X2744 5595 5527 2 1 5467 5176 MUX2 $T=943640 1011480 1 180 $X=939300 $Y=1011100
X2745 1019 5442 2 1 5599 5575 MUX2 $T=939920 1061880 0 0 $X=939920 $Y=1061500
X2746 5608 1018 2 1 5547 1012 MUX2 $T=945500 910680 0 180 $X=941160 $Y=905260
X2747 5604 5527 2 1 5563 5500 MUX2 $T=945500 1011480 0 180 $X=941160 $Y=1006060
X2748 5584 991 2 1 5617 1026 MUX2 $T=941160 1082040 0 0 $X=941160 $Y=1081660
X2749 5613 5609 2 1 5593 5594 MUX2 $T=947360 940920 0 180 $X=943020 $Y=935500
X2750 5597 5457 2 1 5619 5618 MUX2 $T=943640 961080 1 0 $X=943640 $Y=955660
X2751 5596 5562 2 1 5570 5598 MUX2 $T=947980 1021560 0 180 $X=943640 $Y=1016140
X2752 5633 5627 2 1 5557 5395 MUX2 $T=947980 1041720 1 180 $X=943640 $Y=1041340
X2753 5622 5627 2 1 5648 970 MUX2 $T=947360 1031640 0 0 $X=947360 $Y=1031260
X2754 5664 1029 2 1 5624 1012 MUX2 $T=953560 900600 1 180 $X=949220 $Y=900220
X2755 5667 5603 2 1 5645 5618 MUX2 $T=954800 951000 1 180 $X=950460 $Y=950620
X2756 5536 5678 2 1 5628 5258 MUX2 $T=956660 971160 1 180 $X=952320 $Y=970780
X2757 5659 5657 2 1 5680 5395 MUX2 $T=952320 1051800 1 0 $X=952320 $Y=1046380
X2758 5676 1036 2 1 5630 841 MUX2 $T=956660 1082040 0 180 $X=952320 $Y=1076620
X2759 5662 5562 2 1 5679 5500 MUX2 $T=952940 1011480 1 0 $X=952940 $Y=1006060
X2760 5665 5635 2 1 5700 5618 MUX2 $T=954180 940920 1 0 $X=954180 $Y=935500
X2761 5653 5610 2 1 5666 5618 MUX2 $T=958520 961080 0 180 $X=954180 $Y=955660
X2762 5671 5669 2 1 5689 5618 MUX2 $T=956040 920760 0 0 $X=956040 $Y=920380
X2763 1043 5657 2 1 5675 5575 MUX2 $T=960380 1061880 1 180 $X=956040 $Y=1061500
X2764 1039 5657 2 1 5579 970 MUX2 $T=956660 1041720 1 0 $X=956660 $Y=1036300
X2765 5726 5669 2 1 5705 5498 MUX2 $T=965960 920760 1 180 $X=961620 $Y=920380
X2766 1047 1050 2 1 1057 5718 MUX2 $T=962240 1082040 1 0 $X=962240 $Y=1076620
X2767 1048 5635 2 1 5740 5498 MUX2 $T=962860 940920 1 0 $X=962860 $Y=935500
X2768 5727 5610 2 1 5748 5498 MUX2 $T=965340 951000 1 0 $X=965340 $Y=945580
X2769 1063 5721 2 1 5694 5729 MUX2 $T=969680 971160 1 180 $X=965340 $Y=970780
X2770 5731 1036 2 1 5747 5746 MUX2 $T=965340 1071960 1 0 $X=965340 $Y=1066540
X2771 5733 5721 2 1 5754 5598 MUX2 $T=965960 1011480 0 0 $X=965960 $Y=1011100
X2772 1062 5669 2 1 5770 5594 MUX2 $T=969680 930840 1 0 $X=969680 $Y=925420
X2773 5749 5610 2 1 5766 5594 MUX2 $T=970300 951000 1 0 $X=970300 $Y=945580
X2774 5750 5603 2 1 5760 5594 MUX2 $T=970300 951000 0 0 $X=970300 $Y=950620
X2775 5723 1050 2 1 5773 5746 MUX2 $T=970300 1071960 1 0 $X=970300 $Y=1066540
X2776 5759 5657 2 1 5772 5777 MUX2 $T=971540 1051800 1 0 $X=971540 $Y=1046380
X2777 5761 5657 2 1 5781 971 MUX2 $T=972160 1041720 1 0 $X=972160 $Y=1036300
X2778 5788 5779 2 1 5738 5598 MUX2 $T=978360 1011480 1 180 $X=974020 $Y=1011100
X2779 5774 1029 2 1 5792 1072 MUX2 $T=975260 910680 0 0 $X=975260 $Y=910300
X2780 1070 5627 2 1 5806 5777 MUX2 $T=975880 1051800 1 0 $X=975880 $Y=1046380
X2781 5782 5627 2 1 5798 5746 MUX2 $T=975880 1071960 1 0 $X=975880 $Y=1066540
X2782 5795 5796 2 1 5783 5598 MUX2 $T=980840 1001400 1 180 $X=976500 $Y=1001020
X2783 5801 5796 2 1 5811 5729 MUX2 $T=980840 981240 1 0 $X=980840 $Y=975820
X2784 5827 1077 2 1 5803 1072 MUX2 $T=988280 910680 0 180 $X=983940 $Y=905260
X2785 5840 5829 2 1 5832 5729 MUX2 $T=991380 1031640 1 0 $X=991380 $Y=1026220
X2786 5864 5867 2 1 5800 5718 MUX2 $T=996340 1082040 0 180 $X=992000 $Y=1076620
X2787 5894 1084 2 1 5799 5809 MUX2 $T=997580 1061880 1 180 $X=993240 $Y=1061500
X2788 5818 5857 2 1 5849 5729 MUX2 $T=999440 1021560 0 180 $X=995100 $Y=1016140
X2789 5845 1084 2 1 5882 5777 MUX2 $T=995100 1041720 0 0 $X=995100 $Y=1041340
X2790 5888 5867 2 1 5816 1059 MUX2 $T=1000680 1071960 1 180 $X=996340 $Y=1071580
X2791 5895 5867 2 1 5859 5809 MUX2 $T=1001920 1061880 0 180 $X=997580 $Y=1056460
X2792 1096 5867 2 1 5812 5777 MUX2 $T=1003160 1051800 0 180 $X=998820 $Y=1046380
X2793 5917 5921 2 1 5826 1072 MUX2 $T=1005020 920760 0 180 $X=1000680 $Y=915340
X2794 5913 1108 2 1 5881 5900 MUX2 $T=1006880 1031640 0 180 $X=1002540 $Y=1026220
X2795 5945 1084 2 1 5955 1121 MUX2 $T=1007500 1082040 1 0 $X=1007500 $Y=1076620
X2796 5953 5897 2 1 5979 5976 MUX2 $T=1009980 1041720 1 0 $X=1009980 $Y=1036300
X2797 1122 5867 2 1 5989 1130 MUX2 $T=1011220 1082040 0 0 $X=1011220 $Y=1081660
X2798 1124 5867 2 1 5993 1121 MUX2 $T=1012460 1082040 1 0 $X=1012460 $Y=1076620
X2799 6005 1129 2 1 5951 5976 MUX2 $T=1018660 1041720 1 180 $X=1014320 $Y=1041340
X2800 6011 5986 2 1 5950 5900 MUX2 $T=1019280 1021560 0 180 $X=1014940 $Y=1016140
X2801 5998 1129 2 1 6001 5809 MUX2 $T=1016800 1061880 0 0 $X=1016800 $Y=1061500
X2802 6051 1151 2 1 6034 5976 MUX2 $T=1027960 1041720 1 180 $X=1023620 $Y=1041340
X2803 6061 6027 2 1 6037 5900 MUX2 $T=1029820 1021560 0 180 $X=1025480 $Y=1016140
X2804 6086 6080 2 1 6065 6064 MUX2 $T=1034780 991320 0 180 $X=1030440 $Y=985900
X2805 6095 6080 2 1 6066 5900 MUX2 $T=1034780 1021560 0 180 $X=1030440 $Y=1016140
X2806 6069 1156 2 1 6090 5976 MUX2 $T=1031060 1041720 0 0 $X=1031060 $Y=1041340
X2807 5972 1154 2 1 6054 6099 MUX2 $T=1032920 920760 1 0 $X=1032920 $Y=915340
X2808 6016 1160 2 1 6062 5976 MUX2 $T=1038500 1051800 0 180 $X=1034160 $Y=1046380
X2809 6102 1156 2 1 6120 6097 MUX2 $T=1036640 1061880 0 0 $X=1036640 $Y=1061500
X2810 6110 1163 2 1 6129 6099 MUX2 $T=1038500 920760 1 0 $X=1038500 $Y=915340
X2811 6136 6116 2 1 6114 6064 MUX2 $T=1043460 1001400 1 180 $X=1039120 $Y=1001020
X2812 6109 1169 2 1 6147 970 MUX2 $T=1041600 1041720 0 0 $X=1041600 $Y=1041340
X2813 6155 6142 2 1 6131 6064 MUX2 $T=1047180 1001400 0 180 $X=1042840 $Y=995980
X2814 6137 1169 2 1 6156 1176 MUX2 $T=1043460 1051800 1 0 $X=1043460 $Y=1046380
X2815 1183 6158 2 1 6154 5900 MUX2 $T=1050900 1021560 1 180 $X=1046560 $Y=1021180
X2816 6180 6181 2 1 6160 6099 MUX2 $T=1054000 951000 1 180 $X=1049660 $Y=950620
X2817 6164 1160 2 1 6182 6097 MUX2 $T=1049660 1061880 0 0 $X=1049660 $Y=1061500
X2818 6189 6186 2 1 6115 6099 MUX2 $T=1056480 930840 0 180 $X=1052140 $Y=925420
X2819 6193 6190 2 1 6161 6099 MUX2 $T=1056480 971160 1 180 $X=1052140 $Y=970780
X2820 6204 6202 2 1 6178 6064 MUX2 $T=1059580 991320 0 180 $X=1055240 $Y=985900
X2821 1195 1169 2 1 6179 6097 MUX2 $T=1059580 1071960 0 180 $X=1055240 $Y=1066540
X2822 1191 6197 2 1 6216 6099 MUX2 $T=1055860 920760 0 0 $X=1055860 $Y=920380
X2823 6234 6202 2 1 6176 1192 MUX2 $T=1060200 1051800 1 180 $X=1055860 $Y=1051420
X2824 6218 1188 2 1 6195 1194 MUX2 $T=1062060 900600 1 180 $X=1057720 $Y=900220
X2825 6238 6241 2 1 6208 6064 MUX2 $T=1063920 1001400 0 180 $X=1059580 $Y=995980
X2826 1207 6241 2 1 6215 1192 MUX2 $T=1065160 1051800 0 180 $X=1060820 $Y=1046380
X2827 6256 6240 2 1 6222 1176 MUX2 $T=1067020 1011480 1 180 $X=1062680 $Y=1011100
X2828 6239 6240 2 1 6263 6227 MUX2 $T=1063920 1031640 0 0 $X=1063920 $Y=1031260
X2829 6266 6265 2 1 6242 1192 MUX2 $T=1068260 1071960 0 180 $X=1063920 $Y=1066540
X2830 6250 6240 2 1 6273 5777 MUX2 $T=1065160 1051800 1 0 $X=1065160 $Y=1046380
X2831 6274 1210 2 1 6254 1194 MUX2 $T=1070740 900600 1 180 $X=1066400 $Y=900220
X2832 6282 6265 2 1 6247 6097 MUX2 $T=1073220 1071960 0 180 $X=1068880 $Y=1066540
X2833 6253 6265 2 1 6276 5777 MUX2 $T=1074460 1051800 0 180 $X=1070120 $Y=1046380
X2834 6283 6265 2 1 6297 1221 MUX2 $T=1073220 1071960 1 0 $X=1073220 $Y=1066540
X2835 6317 6240 2 1 1218 1217 MUX2 $T=1081280 1082040 0 180 $X=1076940 $Y=1076620
X2836 6329 6240 2 1 6302 1221 MUX2 $T=1082520 1061880 1 180 $X=1078180 $Y=1061500
X2837 6309 1230 2 1 6310 6330 MUX2 $T=1086860 1021560 0 180 $X=1082520 $Y=1016140
X2838 6345 6168 2 1 6362 6366 MUX2 $T=1086240 951000 1 0 $X=1086240 $Y=945580
X2839 6347 1230 2 1 6365 6227 MUX2 $T=1086240 1041720 1 0 $X=1086240 $Y=1036300
X2840 6364 6240 2 1 6324 6097 MUX2 $T=1090580 1071960 1 180 $X=1086240 $Y=1071580
X2841 6383 6303 2 1 6367 6366 MUX2 $T=1094920 951000 0 180 $X=1090580 $Y=945580
X2842 6387 1245 2 1 6340 1239 MUX2 $T=1094920 1071960 1 180 $X=1090580 $Y=1071580
X2843 6385 1234 2 1 6353 6227 MUX2 $T=1095540 1041720 0 180 $X=1091200 $Y=1036300
X2844 1240 6241 2 1 6394 1239 MUX2 $T=1091820 1061880 0 0 $X=1091820 $Y=1061500
X2845 1251 1193 2 1 6355 1244 MUX2 $T=1098640 900600 1 180 $X=1094300 $Y=900220
X2846 6357 1245 2 1 6428 6227 MUX2 $T=1095540 1041720 1 0 $X=1095540 $Y=1036300
X2847 1264 6441 2 1 6417 1239 MUX2 $T=1104220 1061880 1 180 $X=1099880 $Y=1061500
X2848 6423 1245 2 1 6445 1266 MUX2 $T=1101740 1082040 1 0 $X=1101740 $Y=1076620
X2849 1269 1267 2 1 6358 1244 MUX2 $T=1106700 900600 1 180 $X=1102360 $Y=900220
X2850 6432 6370 2 1 6455 1265 MUX2 $T=1103600 930840 0 0 $X=1103600 $Y=930460
X2851 6437 1245 2 1 6456 6330 MUX2 $T=1104220 1021560 1 0 $X=1104220 $Y=1016140
X2852 6464 1193 2 1 6438 1265 MUX2 $T=1109180 920760 0 180 $X=1104840 $Y=915340
X2853 6443 6441 2 1 6458 5821 MUX2 $T=1104840 1051800 1 0 $X=1104840 $Y=1046380
X2854 6459 1268 2 1 6392 1266 MUX2 $T=1109180 1071960 0 180 $X=1104840 $Y=1066540
X2855 6444 1268 2 1 6465 6442 MUX2 $T=1105460 1031640 0 0 $X=1105460 $Y=1031260
X2856 6466 1234 2 1 1277 1238 MUX2 $T=1109180 1082040 0 0 $X=1109180 $Y=1081660
X2857 6475 6359 2 1 6497 1265 MUX2 $T=1111040 930840 1 0 $X=1111040 $Y=925420
X2858 6473 6441 2 1 6499 1238 MUX2 $T=1111040 1051800 0 0 $X=1111040 $Y=1051420
X2859 6476 6241 2 1 6498 1238 MUX2 $T=1111040 1061880 0 0 $X=1111040 $Y=1061500
X2860 6483 6241 2 1 6503 5821 MUX2 $T=1112280 1051800 1 0 $X=1112280 $Y=1046380
X2861 6484 1245 2 1 6504 1238 MUX2 $T=1112280 1071960 1 0 $X=1112280 $Y=1066540
X2862 6493 6441 2 1 6514 6442 MUX2 $T=1114140 1041720 1 0 $X=1114140 $Y=1036300
X2863 1280 1267 2 1 6515 1279 MUX2 $T=1116000 900600 0 0 $X=1116000 $Y=900220
X2864 6406 6486 2 1 6517 6330 MUX2 $T=1116620 1011480 0 0 $X=1116620 $Y=1011100
X2865 6518 6441 2 1 6524 6330 MUX2 $T=1120960 1011480 0 0 $X=1120960 $Y=1011100
X2866 6516 1267 2 1 6527 1265 MUX2 $T=1122820 910680 0 0 $X=1122820 $Y=910300
X2867 6520 6510 2 1 6528 6366 MUX2 $T=1125300 940920 0 0 $X=1125300 $Y=940540
X2868 6525 6255 2 1 6530 6366 MUX2 $T=1125300 951000 0 0 $X=1125300 $Y=950620
X2869 14 11 1364 1403 1 1378 2 AOI22S $T=233120 1041720 1 0 $X=233120 $Y=1036300
X2870 29 1538 1513 1544 1 1417 2 AOI22S $T=254200 1031640 1 0 $X=254200 $Y=1026220
X2871 40 34 1579 1403 1 1378 2 AOI22S $T=263500 1031640 1 180 $X=259780 $Y=1031260
X2872 41 40 1602 1541 1 1609 2 AOI22S $T=263500 1021560 1 0 $X=263500 $Y=1016140
X2873 1604 1617 1542 1619 1 44 2 AOI22S $T=265360 920760 1 0 $X=265360 $Y=915340
X2874 1576 1615 1610 43 1 53 2 AOI22S $T=267220 951000 0 0 $X=267220 $Y=950620
X2875 1452 1677 1726 1717 1 1586 2 AOI22S $T=283960 1041720 1 180 $X=280240 $Y=1041340
X2876 1779 1774 1783 1814 1 1792 2 AOI22S $T=290780 1051800 0 0 $X=290780 $Y=1051420
X2877 1803 1811 1683 1856 1 1819 2 AOI22S $T=293880 961080 0 0 $X=293880 $Y=960700
X2878 1792 1821 1814 1827 1 1779 2 AOI22S $T=295120 1041720 0 0 $X=295120 $Y=1041340
X2879 1820 46 1831 1796 1 1674 2 AOI22S $T=298220 1031640 1 0 $X=298220 $Y=1026220
X2880 1894 1872 1833 1866 1 1714 2 AOI22S $T=305660 940920 0 180 $X=301940 $Y=935500
X2881 1876 1883 1812 1777 1 1861 2 AOI22S $T=303800 971160 1 0 $X=303800 $Y=965740
X2882 90 94 1646 1906 1 98 2 AOI22S $T=309380 930840 1 0 $X=309380 $Y=925420
X2883 101 1902 1818 105 1 90 2 AOI22S $T=312480 930840 0 0 $X=312480 $Y=930460
X2884 1902 90 1757 1943 1 94 2 AOI22S $T=312480 951000 1 0 $X=312480 $Y=945580
X2885 1749 79 1901 1913 1 1808 2 AOI22S $T=314340 1031640 1 0 $X=314340 $Y=1026220
X2886 1749 79 1998 1800 1 1912 2 AOI22S $T=324880 1031640 0 180 $X=321160 $Y=1026220
X2887 1986 2014 2039 2000 1 1985 2 AOI22S $T=332320 940920 0 180 $X=328600 $Y=935500
X2888 145 155 156 2135 1 2137 2 AOI22S $T=345960 1082040 1 180 $X=342240 $Y=1081660
X2889 119 129 2161 1912 1 1913 2 AOI22S $T=347200 1031640 0 180 $X=343480 $Y=1026220
X2890 2200 2212 2153 2209 1 2188 2 AOI22S $T=357740 951000 0 180 $X=354020 $Y=945580
X2891 2262 2213 2240 178 1 2229 2 AOI22S $T=365180 951000 1 180 $X=361460 $Y=950620
X2892 2269 2276 2282 2265 1 2238 2 AOI22S $T=367040 940920 0 0 $X=367040 $Y=940540
X2893 2228 2322 2353 2351 1 2363 2 AOI22S $T=376960 940920 1 0 $X=376960 $Y=935500
X2894 2433 2419 2435 2406 1 2374 2 AOI22S $T=392460 1041720 1 180 $X=388740 $Y=1041340
X2895 2446 208 2436 2330 1 2329 2 AOI22S $T=392460 1071960 1 180 $X=388740 $Y=1071580
X2896 2433 2419 2466 2457 1 2349 2 AOI22S $T=396180 1041720 1 180 $X=392460 $Y=1041340
X2897 2433 2419 2482 2348 1 2243 2 AOI22S $T=399900 1041720 1 180 $X=396180 $Y=1041340
X2898 2539 2523 225 2520 1 2256 2 AOI22S $T=407340 1011480 0 180 $X=403620 $Y=1006060
X2899 2539 2523 2554 2534 1 2461 2 AOI22S $T=411060 1011480 1 180 $X=407340 $Y=1011100
X2900 2579 2561 2566 2498 1 2452 2 AOI22S $T=412920 981240 0 180 $X=409200 $Y=975820
X2901 2540 2523 2574 2551 1 2501 2 AOI22S $T=414160 1001400 1 180 $X=410440 $Y=1001020
X2902 2539 2523 2560 2526 1 2300 2 AOI22S $T=414160 1041720 0 180 $X=410440 $Y=1036300
X2903 2433 2556 232 2541 1 2313 2 AOI22S $T=414780 1051800 0 180 $X=411060 $Y=1046380
X2904 2579 2561 2581 2477 1 2290 2 AOI22S $T=413540 981240 1 0 $X=413540 $Y=975820
X2905 2579 2561 2643 2638 1 2458 2 AOI22S $T=424700 971160 1 180 $X=420980 $Y=970780
X2906 2680 2556 2714 2658 1 2493 2 AOI22S $T=436480 1031640 1 180 $X=432760 $Y=1031260
X2907 2680 2721 2716 2694 1 2705 2 AOI22S $T=435240 1031640 1 0 $X=435240 $Y=1026220
X2908 2728 254 2724 258 1 242 2 AOI22S $T=438960 1071960 1 180 $X=435240 $Y=1071580
X2909 2710 2721 2737 2729 1 2382 2 AOI22S $T=440820 991320 1 180 $X=437100 $Y=990940
X2910 2767 2561 2770 2662 1 2612 2 AOI22S $T=446400 961080 0 180 $X=442680 $Y=955660
X2911 2767 2768 2775 2704 1 2743 2 AOI22S $T=447640 971160 1 180 $X=443920 $Y=970780
X2912 2680 2556 2761 2689 1 2274 2 AOI22S $T=443920 1031640 0 0 $X=443920 $Y=1031260
X2913 2728 2483 2763 2589 1 271 2 AOI22S $T=444540 1071960 0 0 $X=444540 $Y=1071580
X2914 2767 2561 2802 2774 1 2722 2 AOI22S $T=451360 961080 0 180 $X=447640 $Y=955660
X2915 2710 2721 2815 2795 1 2757 2 AOI22S $T=452600 991320 1 180 $X=448880 $Y=990940
X2916 2540 273 2801 2703 1 2817 2 AOI22S $T=451360 940920 0 0 $X=451360 $Y=940540
X2917 2767 2561 2824 2438 1 2833 2 AOI22S $T=454460 961080 1 0 $X=454460 $Y=955660
X2918 2540 273 2826 2410 1 2532 2 AOI22S $T=455080 940920 0 0 $X=455080 $Y=940540
X2919 289 286 2866 2726 1 2687 2 AOI22S $T=464380 920760 0 180 $X=460660 $Y=915340
X2920 289 286 2874 275 1 2742 2 AOI22S $T=465620 920760 1 180 $X=461900 $Y=920380
X2921 2908 2884 2891 2830 1 2889 2 AOI22S $T=472440 991320 0 180 $X=468720 $Y=985900
X2922 2908 2884 2927 2911 1 2880 2 AOI22S $T=473680 1001400 1 180 $X=469960 $Y=1001020
X2923 2908 2904 2913 2907 1 2933 2 AOI22S $T=471820 1031640 1 0 $X=471820 $Y=1026220
X2924 2984 311 2978 2965 1 2916 2 AOI22S $T=483600 940920 1 180 $X=479880 $Y=940540
X2925 312 313 2919 2975 1 2974 2 AOI22S $T=485460 920760 1 180 $X=481740 $Y=920380
X2926 2710 2979 2896 2985 1 2989 2 AOI22S $T=482360 1011480 0 0 $X=482360 $Y=1011100
X2927 312 313 2924 2660 1 317 2 AOI22S $T=482980 910680 0 0 $X=482980 $Y=910300
X2928 2710 2721 2995 3020 1 2963 2 AOI22S $T=485460 991320 1 0 $X=485460 $Y=985900
X2929 2984 311 3007 3013 1 3021 2 AOI22S $T=488560 951000 1 0 $X=488560 $Y=945580
X2930 2579 2884 3019 2959 1 2994 2 AOI22S $T=490420 981240 1 0 $X=490420 $Y=975820
X2931 289 2884 333 3099 1 2584 2 AOI22S $T=503440 920760 0 0 $X=503440 $Y=920380
X2932 343 340 344 3112 1 330 2 AOI22S $T=507160 910680 0 0 $X=507160 $Y=910300
X2933 3182 3166 3173 358 1 3117 2 AOI22S $T=520800 1001400 0 180 $X=517080 $Y=995980
X2934 3185 3177 3155 3174 1 3153 2 AOI22S $T=522660 1051800 1 180 $X=518940 $Y=1051420
X2935 3185 3177 3163 3160 1 337 2 AOI22S $T=523280 1071960 0 180 $X=519560 $Y=1066540
X2936 3182 3166 3205 3143 1 3151 2 AOI22S $T=524520 1001400 0 180 $X=520800 $Y=995980
X2937 3185 3177 3197 3207 1 3125 2 AOI22S $T=523280 1071960 0 0 $X=523280 $Y=1071580
X2938 3182 3166 3216 2509 1 2413 2 AOI22S $T=527620 971160 1 180 $X=523900 $Y=970780
X2939 3185 3192 3208 3171 1 3189 2 AOI22S $T=524520 1041720 1 0 $X=524520 $Y=1036300
X2940 3182 3166 3227 2189 1 366 2 AOI22S $T=530720 981240 1 180 $X=527000 $Y=980860
X2941 343 340 369 3178 1 3212 2 AOI22S $T=528860 910680 1 0 $X=528860 $Y=905260
X2942 3203 3233 3237 3156 1 3188 2 AOI22S $T=533820 951000 0 180 $X=530100 $Y=945580
X2943 3203 3233 3238 3183 1 2365 2 AOI22S $T=534440 940920 1 180 $X=530720 $Y=940540
X2944 3182 3233 3239 3214 1 2272 2 AOI22S $T=534440 971160 1 180 $X=530720 $Y=970780
X2945 3182 3166 3244 3236 1 3199 2 AOI22S $T=534440 981240 1 180 $X=530720 $Y=980860
X2946 3203 3233 3226 2123 1 2261 2 AOI22S $T=531340 951000 0 0 $X=531340 $Y=950620
X2947 387 384 3268 382 1 3250 2 AOI22S $T=538780 1071960 1 180 $X=535060 $Y=1071580
X2948 3291 3283 3242 390 1 378 2 AOI22S $T=542500 1011480 1 180 $X=538780 $Y=1011100
X2949 3311 3293 3234 2219 1 3284 2 AOI22S $T=544360 1001400 0 180 $X=540640 $Y=995980
X2950 3271 3192 3304 3269 1 3235 2 AOI22S $T=544980 1051800 0 180 $X=541260 $Y=1046380
X2951 3291 3283 3326 408 1 2236 2 AOI22S $T=546840 1011480 0 0 $X=546840 $Y=1011100
X2952 415 403 3341 3299 1 3330 2 AOI22S $T=551180 940920 1 180 $X=547460 $Y=940540
X2953 407 3336 3289 3315 1 2305 2 AOI22S $T=551180 971160 1 180 $X=547460 $Y=970780
X2954 3311 3293 3331 3308 1 2231 2 AOI22S $T=551180 1001400 1 0 $X=551180 $Y=995980
X2955 3377 3293 3310 3365 1 3329 2 AOI22S $T=557380 940920 1 180 $X=553660 $Y=940540
X2956 332 403 3418 421 1 419 2 AOI22S $T=561100 900600 1 180 $X=557380 $Y=900220
X2957 3364 413 3384 3390 1 2674 2 AOI22S $T=558000 961080 1 0 $X=558000 $Y=955660
X2958 3396 3192 3388 3371 1 3412 2 AOI22S $T=559240 1061880 1 0 $X=559240 $Y=1056460
X2959 3396 3192 3386 3416 1 3410 2 AOI22S $T=562960 1051800 0 0 $X=562960 $Y=1051420
X2960 3291 3283 3426 3434 1 3423 2 AOI22S $T=564200 1011480 0 0 $X=564200 $Y=1011100
X2961 3396 3400 3429 3357 1 425 2 AOI22S $T=567920 1071960 1 180 $X=564200 $Y=1071580
X2962 3291 3283 3445 3344 1 429 2 AOI22S $T=568540 1021560 1 180 $X=564820 $Y=1021180
X2963 3377 3293 3393 2598 1 435 2 AOI22S $T=565440 951000 1 0 $X=565440 $Y=945580
X2964 387 384 3436 3322 1 3448 2 AOI22S $T=566060 1082040 1 0 $X=566060 $Y=1076620
X2965 407 3437 3455 3408 1 437 2 AOI22S $T=571640 981240 0 180 $X=567920 $Y=975820
X2966 3291 3283 3454 436 1 440 2 AOI22S $T=569160 1021560 0 0 $X=569160 $Y=1021180
X2967 415 403 3456 3435 1 3466 2 AOI22S $T=569780 920760 1 0 $X=569780 $Y=915340
X2968 3443 3437 3477 445 1 446 2 AOI22S $T=573500 1001400 1 0 $X=573500 $Y=995980
X2969 3377 3293 3459 3478 1 3218 2 AOI22S $T=574120 951000 1 0 $X=574120 $Y=945580
X2970 3396 3400 442 450 1 448 2 AOI22S $T=574120 1082040 1 0 $X=574120 $Y=1076620
X2971 3443 3437 3480 3468 1 3490 2 AOI22S $T=574740 991320 1 0 $X=574740 $Y=985900
X2972 3443 3437 3482 3481 1 452 2 AOI22S $T=575980 971160 0 0 $X=575980 $Y=970780
X2973 3271 3500 3494 3499 1 3510 2 AOI22S $T=579700 1021560 1 0 $X=579700 $Y=1016140
X2974 3271 3400 3483 3524 1 3534 2 AOI22S $T=580320 1021560 0 0 $X=580320 $Y=1021180
X2975 3377 3519 3484 3514 1 2496 2 AOI22S $T=582800 961080 1 0 $X=582800 $Y=955660
X2976 3396 3400 3512 438 1 3507 2 AOI22S $T=582800 1061880 1 0 $X=582800 $Y=1056460
X2977 3532 3500 3430 3544 1 476 2 AOI22S $T=585900 981240 0 0 $X=585900 $Y=980860
X2978 473 469 3518 3462 1 2631 2 AOI22S $T=586520 920760 1 0 $X=586520 $Y=915340
X2979 473 469 3541 3529 1 478 2 AOI22S $T=587140 930840 0 0 $X=587140 $Y=930460
X2980 473 469 475 477 1 479 2 AOI22S $T=587760 900600 0 0 $X=587760 $Y=900220
X2981 3532 3519 3476 3546 1 471 2 AOI22S $T=588380 971160 1 0 $X=588380 $Y=965740
X2982 3532 3500 3497 3552 1 481 2 AOI22S $T=589620 981240 0 0 $X=589620 $Y=980860
X2983 484 413 3528 2597 1 3603 2 AOI22S $T=598920 920760 1 0 $X=598920 $Y=915340
X2984 484 413 3503 3621 1 3627 2 AOI22S $T=603880 910680 1 0 $X=603880 $Y=905260
X2985 3674 3656 3664 3641 1 3619 2 AOI22S $T=613800 1051800 0 180 $X=610080 $Y=1046380
X2986 3674 3656 3700 3571 1 508 2 AOI22S $T=618140 1051800 0 180 $X=614420 $Y=1046380
X2987 3696 3706 3709 3660 1 3588 2 AOI22S $T=620620 1041720 0 180 $X=616900 $Y=1036300
X2988 3696 3706 3699 3670 1 3611 2 AOI22S $T=617520 1031640 0 0 $X=617520 $Y=1031260
X2989 3754 3741 3761 505 1 3692 2 AOI22S $T=626200 971160 1 180 $X=622480 $Y=970780
X2990 3754 3741 3773 3724 1 3487 2 AOI22S $T=629300 961080 1 180 $X=625580 $Y=960700
X2991 3774 3757 3745 3550 1 510 2 AOI22S $T=629300 1011480 0 180 $X=625580 $Y=1006060
X2992 3696 3706 3718 3738 1 3764 2 AOI22S $T=625580 1041720 1 0 $X=625580 $Y=1036300
X2993 3778 3765 3756 3728 1 3691 2 AOI22S $T=630540 951000 0 180 $X=626820 $Y=945580
X2994 3774 3757 3781 521 1 511 2 AOI22S $T=633020 1011480 0 180 $X=629300 $Y=1006060
X2995 3696 3706 3737 537 1 535 2 AOI22S $T=629300 1031640 0 0 $X=629300 $Y=1031260
X2996 3778 3765 3788 525 1 539 2 AOI22S $T=634260 951000 1 180 $X=630540 $Y=950620
X2997 3778 3765 3799 531 1 3785 2 AOI22S $T=635500 951000 0 180 $X=631780 $Y=945580
X2998 3758 3748 3783 3694 1 3569 2 AOI22S $T=631780 991320 1 0 $X=631780 $Y=985900
X2999 3774 3757 3802 3790 1 3766 2 AOI22S $T=638600 1011480 0 180 $X=634880 $Y=1006060
X3000 3758 3748 3796 550 1 553 2 AOI22S $T=635500 991320 1 0 $X=635500 $Y=985900
X3001 3754 3741 3814 552 1 555 2 AOI22S $T=642940 971160 1 180 $X=639220 $Y=970780
X3002 3836 3832 3843 3771 1 3791 2 AOI22S $T=645420 1051800 1 180 $X=641700 $Y=1051420
X3003 574 572 3868 570 1 3776 2 AOI22S $T=652860 920760 0 180 $X=649140 $Y=915340
X3004 3754 3741 3882 3599 1 3869 2 AOI22S $T=655340 971160 0 180 $X=651620 $Y=965740
X3005 574 572 578 3848 1 563 2 AOI22S $T=655960 900600 1 180 $X=652240 $Y=900220
X3006 3841 3706 3888 3880 1 3596 2 AOI22S $T=655960 1031640 1 180 $X=652240 $Y=1031260
X3007 3758 3748 3879 3607 1 3733 2 AOI22S $T=652860 991320 1 0 $X=652860 $Y=985900
X3008 3774 3757 3892 3884 1 581 2 AOI22S $T=654720 1011480 1 0 $X=654720 $Y=1006060
X3009 574 572 3921 3902 1 579 2 AOI22S $T=659680 900600 1 180 $X=655960 $Y=900220
X3010 587 585 3913 3573 1 3643 2 AOI22S $T=660300 940920 0 180 $X=656580 $Y=935500
X3011 3754 3741 3910 3873 1 3922 2 AOI22S $T=657820 971160 1 0 $X=657820 $Y=965740
X3012 3774 3757 3928 3639 1 3934 2 AOI22S $T=660300 1011480 1 0 $X=660300 $Y=1006060
X3013 3778 585 3932 3883 1 564 2 AOI22S $T=662160 951000 1 0 $X=662160 $Y=945580
X3014 3758 3748 3930 3563 1 592 2 AOI22S $T=662160 981240 0 0 $X=662160 $Y=980860
X3015 3841 3947 3948 3978 1 3918 2 AOI22S $T=664640 1041720 1 0 $X=664640 $Y=1036300
X3016 4011 4005 611 3937 1 4001 2 AOI22S $T=675180 971160 0 180 $X=671460 $Y=965740
X3017 4020 4005 615 3970 1 4001 2 AOI22S $T=676420 961080 0 180 $X=672700 $Y=955660
X3018 4023 3991 617 4005 1 4001 2 AOI22S $T=677040 961080 1 180 $X=673320 $Y=960700
X3019 4049 4005 625 3989 1 4001 2 AOI22S $T=680760 951000 1 180 $X=677040 $Y=950620
X3020 4029 4008 4038 4043 1 4000 2 AOI22S $T=682000 991320 0 180 $X=678280 $Y=985900
X3021 626 601 4067 3945 1 3982 2 AOI22S $T=683860 920760 0 180 $X=680140 $Y=915340
X3022 3891 601 4028 628 1 4063 2 AOI22S $T=680140 971160 1 0 $X=680140 $Y=965740
X3023 3999 3961 4031 3898 1 3609 2 AOI22S $T=680760 951000 0 0 $X=680760 $Y=950620
X3024 3841 3947 4057 4040 1 640 2 AOI22S $T=681380 1041720 1 0 $X=681380 $Y=1036300
X3025 3836 3832 4065 632 1 618 2 AOI22S $T=682620 1051800 1 0 $X=682620 $Y=1046380
X3026 3891 601 4070 3993 1 4095 2 AOI22S $T=684480 951000 0 0 $X=684480 $Y=950620
X3027 3774 3757 4083 639 1 3808 2 AOI22S $T=685100 1011480 1 0 $X=685100 $Y=1006060
X3028 3841 3947 4098 4085 1 4009 2 AOI22S $T=688820 1031640 0 0 $X=688820 $Y=1031260
X3029 4078 4100 4044 4051 1 3949 2 AOI22S $T=689440 1011480 1 0 $X=689440 $Y=1006060
X3030 3836 3832 4091 4120 1 3992 2 AOI22S $T=690060 1051800 1 0 $X=690060 $Y=1046380
X3031 4029 4008 4082 4127 1 4108 2 AOI22S $T=692540 991320 1 0 $X=692540 $Y=985900
X3032 4159 3947 4170 4178 1 4148 2 AOI22S $T=699980 1041720 1 0 $X=699980 $Y=1036300
X3033 4126 4041 4222 4197 1 4211 2 AOI22S $T=711140 961080 1 180 $X=707420 $Y=960700
X3034 4139 4158 4181 4225 1 4052 2 AOI22S $T=707420 1051800 0 0 $X=707420 $Y=1051420
X3035 662 663 4168 664 1 4147 2 AOI22S $T=708040 910680 1 0 $X=708040 $Y=905260
X3036 662 663 4138 4140 1 3907 2 AOI22S $T=708040 920760 1 0 $X=708040 $Y=915340
X3037 3999 3961 4237 4203 1 4223 2 AOI22S $T=713620 940920 1 180 $X=709900 $Y=940540
X3038 4029 4226 4243 4224 1 665 2 AOI22S $T=713620 981240 1 180 $X=709900 $Y=980860
X3039 4126 4041 4249 4198 1 4235 2 AOI22S $T=715480 971160 1 180 $X=711760 $Y=970780
X3040 4126 4041 4234 666 1 4252 2 AOI22S $T=713000 951000 0 0 $X=713000 $Y=950620
X3041 4078 4100 4242 4238 1 670 2 AOI22S $T=713620 1001400 0 0 $X=713620 $Y=1001020
X3042 662 4226 4284 4233 1 4115 2 AOI22S $T=721680 920760 1 180 $X=717960 $Y=920380
X3043 4278 4271 4275 673 1 4194 2 AOI22S $T=721680 1031640 0 180 $X=717960 $Y=1026220
X3044 4299 676 678 3990 1 4001 2 AOI22S $T=722920 951000 0 180 $X=719200 $Y=945580
X3045 3999 3961 4274 4282 1 4287 2 AOI22S $T=720440 940920 0 0 $X=720440 $Y=940540
X3046 4139 4158 4326 4285 1 681 2 AOI22S $T=725400 1061880 0 180 $X=721680 $Y=1056460
X3047 4139 4158 4289 4333 1 4323 2 AOI22S $T=724780 1031640 0 0 $X=724780 $Y=1031260
X3048 662 4226 4286 4320 1 4305 2 AOI22S $T=725400 981240 1 0 $X=725400 $Y=975820
X3049 4310 4328 689 693 1 691 2 AOI22S $T=727260 910680 1 0 $X=727260 $Y=905260
X3050 4310 4328 4145 4309 1 4335 2 AOI22S $T=727260 920760 1 0 $X=727260 $Y=915340
X3051 4310 4328 4292 4334 1 4266 2 AOI22S $T=727260 991320 1 0 $X=727260 $Y=985900
X3052 4139 4100 4330 4046 1 4343 2 AOI22S $T=727880 1001400 1 0 $X=727880 $Y=995980
X3053 4310 4328 4311 4301 1 4345 2 AOI22S $T=728500 920760 0 0 $X=728500 $Y=920380
X3054 662 4226 4327 3577 1 690 2 AOI22S $T=729120 971160 1 0 $X=729120 $Y=965740
X3055 4278 4271 4348 695 1 4370 2 AOI22S $T=730980 1031640 1 0 $X=730980 $Y=1026220
X3056 702 694 4174 703 1 4394 2 AOI22S $T=735940 910680 1 0 $X=735940 $Y=905260
X3057 4557 4544 4548 730 1 4516 2 AOI22S $T=770660 1031640 1 180 $X=766940 $Y=1031260
X3058 4565 4544 4559 745 1 4483 2 AOI22S $T=770660 1071960 0 180 $X=766940 $Y=1066540
X3059 4555 4543 4551 4456 1 746 2 AOI22S $T=771280 991320 1 180 $X=767560 $Y=990940
X3060 4565 4544 4558 4502 1 744 2 AOI22S $T=771280 1061880 0 180 $X=767560 $Y=1056460
X3061 4555 4540 4561 4448 1 733 2 AOI22S $T=771900 971160 1 180 $X=768180 $Y=970780
X3062 4576 4540 4572 4486 1 751 2 AOI22S $T=773760 951000 1 180 $X=770040 $Y=950620
X3063 754 753 4573 4512 1 714 2 AOI22S $T=773760 1082040 0 180 $X=770040 $Y=1076620
X3064 4576 4540 4586 4525 1 4492 2 AOI22S $T=774380 961080 1 180 $X=770660 $Y=960700
X3065 4555 4543 4574 4012 1 756 2 AOI22S $T=771900 991320 0 0 $X=771900 $Y=990940
X3066 4600 4597 4616 4504 1 760 2 AOI22S $T=778720 930840 1 180 $X=775000 $Y=930460
X3067 4557 4544 4594 4501 1 4585 2 AOI22S $T=775620 1041720 0 0 $X=775620 $Y=1041340
X3068 4557 4544 4602 734 1 4580 2 AOI22S $T=775620 1051800 0 0 $X=775620 $Y=1051420
X3069 4624 4005 766 4613 1 4365 2 AOI22S $T=780580 1001400 1 180 $X=776860 $Y=1001020
X3070 4579 4606 4630 4622 1 4541 2 AOI22S $T=782440 1011480 1 180 $X=778720 $Y=1011100
X3071 4579 4633 770 774 1 4610 2 AOI22S $T=780580 900600 0 0 $X=780580 $Y=900220
X3072 4579 4606 4653 4510 1 4526 2 AOI22S $T=784920 1021560 1 180 $X=781200 $Y=1021180
X3073 4600 4597 4678 4569 1 4654 2 AOI22S $T=789880 940920 0 180 $X=786160 $Y=935500
X3074 789 785 4677 4628 1 778 2 AOI22S $T=791120 910680 1 180 $X=787400 $Y=910300
X3075 4600 4597 4728 802 1 797 2 AOI22S $T=796700 940920 0 180 $X=792980 $Y=935500
X3076 789 785 815 4760 1 813 2 AOI22S $T=802900 910680 1 180 $X=799180 $Y=910300
X3077 4813 4823 4828 4786 1 4769 2 AOI22S $T=810340 951000 1 180 $X=806620 $Y=950620
X3078 4813 4782 4831 4632 1 4517 2 AOI22S $T=810340 961080 1 180 $X=806620 $Y=960700
X3079 822 823 4748 4805 1 826 2 AOI22S $T=809720 1082040 1 0 $X=809720 $Y=1076620
X3080 832 4823 4817 4847 1 4554 2 AOI22S $T=814680 930840 1 180 $X=810960 $Y=930460
X3081 822 823 4740 4860 1 834 2 AOI22S $T=813440 1082040 1 0 $X=813440 $Y=1076620
X3082 789 4883 4820 4863 1 4886 2 AOI22S $T=815920 1021560 1 0 $X=815920 $Y=1016140
X3083 4848 4883 4799 844 1 4904 2 AOI22S $T=819020 1031640 0 0 $X=819020 $Y=1031260
X3084 4848 823 4816 4859 1 4873 2 AOI22S $T=819020 1051800 0 0 $X=819020 $Y=1051420
X3085 4924 4823 4887 846 1 4676 2 AOI22S $T=823980 951000 0 180 $X=820260 $Y=945580
X3086 4848 823 4844 4916 1 852 2 AOI22S $T=822740 1051800 0 0 $X=822740 $Y=1051420
X3087 832 4823 4889 4901 1 4922 2 AOI22S $T=823360 930840 0 0 $X=823360 $Y=930460
X3088 4894 4883 4789 4734 1 4903 2 AOI22S $T=823360 1021560 1 0 $X=823360 $Y=1016140
X3089 4997 4992 4993 4750 1 4974 2 AOI22S $T=841340 961080 1 180 $X=837620 $Y=960700
X3090 4600 4597 4987 5001 1 4649 2 AOI22S $T=839480 940920 0 0 $X=839480 $Y=940540
X3091 4959 4995 5014 858 1 5003 2 AOI22S $T=844440 920760 0 180 $X=840720 $Y=915340
X3092 5065 5055 5059 5036 1 5047 2 AOI22S $T=851260 1061880 1 180 $X=847540 $Y=1061500
X3093 5065 5055 5076 4937 1 5045 2 AOI22S $T=852500 1011480 1 180 $X=848780 $Y=1011100
X3094 4997 4992 5062 4783 1 5074 2 AOI22S $T=850640 961080 0 0 $X=850640 $Y=960700
X3095 5065 5055 5077 5005 1 5069 2 AOI22S $T=854980 1041720 1 180 $X=851260 $Y=1041340
X3096 883 886 5082 885 1 874 2 AOI22S $T=854360 1071960 1 0 $X=854360 $Y=1066540
X3097 5065 5101 5107 5094 1 5072 2 AOI22S $T=859320 1011480 1 180 $X=855600 $Y=1011100
X3098 5065 5055 5112 5068 1 5088 2 AOI22S $T=859320 1041720 0 180 $X=855600 $Y=1036300
X3099 4959 4995 5110 891 1 5078 2 AOI22S $T=860560 910680 1 180 $X=856840 $Y=910300
X3100 883 886 5126 865 1 892 2 AOI22S $T=863040 1082040 1 180 $X=859320 $Y=1081660
X3101 4959 4995 897 888 1 5083 2 AOI22S $T=863660 910680 0 180 $X=859940 $Y=905260
X3102 5147 5124 5148 5137 1 5130 2 AOI22S $T=866140 971160 0 180 $X=862420 $Y=965740
X3103 5065 5101 5142 4953 1 902 2 AOI22S $T=863660 1011480 0 0 $X=863660 $Y=1011100
X3104 4997 4992 5159 5104 1 5091 2 AOI22S $T=868620 951000 0 180 $X=864900 $Y=945580
X3105 5147 5124 5191 5221 1 914 2 AOI22S $T=874820 961080 0 0 $X=874820 $Y=960700
X3106 5264 4633 5250 5192 1 5243 2 AOI22S $T=884120 1021560 1 180 $X=880400 $Y=1021180
X3107 5264 5214 5184 5235 1 922 2 AOI22S $T=884740 1041720 0 180 $X=881020 $Y=1036300
X3108 5248 925 5135 5253 1 927 2 AOI22S $T=882880 1071960 1 0 $X=882880 $Y=1066540
X3109 5264 5214 5304 5309 1 5298 2 AOI22S $T=888460 1051800 0 0 $X=888460 $Y=1051420
X3110 5225 5242 5322 5281 1 5290 2 AOI22S $T=892800 951000 1 180 $X=889080 $Y=950620
X3111 5264 4633 5297 5320 1 5325 2 AOI22S $T=890320 1021560 0 0 $X=890320 $Y=1021180
X3112 5225 5242 5342 5330 1 939 2 AOI22S $T=897140 961080 0 180 $X=893420 $Y=955660
X3113 5315 5338 5343 5268 1 940 2 AOI22S $T=897140 991320 0 180 $X=893420 $Y=985900
X3114 5225 5242 5350 942 1 932 2 AOI22S $T=897760 951000 1 180 $X=894040 $Y=950620
X3115 5225 5242 5356 5345 1 949 2 AOI22S $T=897760 951000 0 0 $X=897760 $Y=950620
X3116 5264 4633 5341 951 1 950 2 AOI22S $T=897760 1021560 0 0 $X=897760 $Y=1021180
X3117 5225 5242 5378 5383 1 957 2 AOI22S $T=901480 961080 1 0 $X=901480 $Y=955660
X3118 5315 5338 5400 5397 1 5375 2 AOI22S $T=907680 971160 1 0 $X=907680 $Y=965740
X3119 5315 5338 5360 5377 1 5393 2 AOI22S $T=908300 971160 0 0 $X=908300 $Y=970780
X3120 5315 5338 5401 966 1 5417 2 AOI22S $T=909540 991320 0 0 $X=909540 $Y=990940
X3121 5315 5338 5416 5413 1 5423 2 AOI22S $T=911400 981240 1 0 $X=911400 $Y=975820
X3122 5465 5453 5459 5427 1 5407 2 AOI22S $T=923800 1061880 0 180 $X=920080 $Y=1056460
X3123 982 984 5466 5412 1 5483 2 AOI22S $T=921320 1082040 1 0 $X=921320 $Y=1076620
X3124 5534 5526 5525 5521 1 5520 2 AOI22S $T=934340 961080 0 180 $X=930620 $Y=955660
X3125 5534 1007 5546 5472 1 5512 2 AOI22S $T=934960 940920 0 180 $X=931240 $Y=935500
X3126 5534 1007 1009 5544 1 1016 2 AOI22S $T=933720 900600 0 0 $X=933720 $Y=900220
X3127 5558 5548 5541 5484 1 1010 2 AOI22S $T=938060 930840 1 180 $X=934340 $Y=930460
X3128 5545 5559 5566 5522 1 5504 2 AOI22S $T=939300 1011480 1 180 $X=935580 $Y=1011100
X3129 5545 5559 5567 990 1 986 2 AOI22S $T=939920 1011480 0 180 $X=936200 $Y=1006060
X3130 5553 5548 5531 5573 1 5569 2 AOI22S $T=936820 940920 0 0 $X=936820 $Y=940540
X3131 5553 5559 5588 5539 1 1014 2 AOI22S $T=941780 991320 0 180 $X=938060 $Y=985900
X3132 5545 5559 5574 5447 1 5488 2 AOI22S $T=938680 1031640 0 0 $X=938680 $Y=1031260
X3133 5534 5526 5591 5582 1 5450 2 AOI22S $T=943640 961080 0 180 $X=939920 $Y=955660
X3134 1000 1007 1025 5612 1 5616 2 AOI22S $T=944880 900600 0 0 $X=944880 $Y=900220
X3135 5654 5526 5606 5629 1 5592 2 AOI22S $T=951080 991320 0 180 $X=947360 $Y=985900
X3136 5654 5646 5611 5638 1 5602 2 AOI22S $T=952320 1011480 0 180 $X=948600 $Y=1006060
X3137 5655 5644 5649 5639 1 5641 2 AOI22S $T=952320 1051800 0 180 $X=948600 $Y=1046380
X3138 5654 5646 5621 5561 1 5529 2 AOI22S $T=952940 1011480 1 180 $X=949220 $Y=1011100
X3139 1021 5548 5642 5631 1 5660 2 AOI22S $T=950460 930840 0 0 $X=950460 $Y=930460
X3140 1028 1031 5661 5677 1 1033 2 AOI22S $T=952320 1071960 0 0 $X=952320 $Y=1071580
X3141 5655 5644 5668 1032 1 5626 2 AOI22S $T=956660 1041720 0 180 $X=952940 $Y=1036300
X3142 5687 5636 5637 5615 1 5672 2 AOI22S $T=959140 951000 1 180 $X=955420 $Y=950620
X3143 1042 1035 1041 1040 1 5681 2 AOI22S $T=960380 900600 1 180 $X=956660 $Y=900220
X3144 5654 5526 5693 5507 1 1046 2 AOI22S $T=959140 971160 0 0 $X=959140 $Y=970780
X3145 1028 1031 5695 5730 1 5699 2 AOI22S $T=959140 1071960 0 0 $X=959140 $Y=1071580
X3146 5654 1031 5706 5685 1 5556 2 AOI22S $T=960380 991320 0 0 $X=960380 $Y=990940
X3147 5655 5644 5709 5722 1 1051 2 AOI22S $T=961000 1041720 0 0 $X=961000 $Y=1041340
X3148 1042 1035 1056 5736 1 5741 2 AOI22S $T=965340 910680 1 0 $X=965340 $Y=905260
X3149 5707 5548 5744 5710 1 1067 2 AOI22S $T=969060 940920 1 0 $X=969060 $Y=935500
X3150 5553 1052 5758 5756 1 5647 2 AOI22S $T=972160 991320 0 0 $X=972160 $Y=990940
X3151 5553 1052 5698 5769 1 5776 2 AOI22S $T=972780 1001400 0 0 $X=972780 $Y=1001020
X3152 5687 5636 5771 5778 1 5786 2 AOI22S $T=974640 951000 0 0 $X=974640 $Y=950620
X3153 5883 5870 5879 5833 1 5813 2 AOI22S $T=1000060 1011480 0 180 $X=996340 $Y=1006060
X3154 5892 5877 1092 1075 1 5842 2 AOI22S $T=1000680 1082040 0 180 $X=996960 $Y=1076620
X3155 5883 5887 5891 5841 1 5808 2 AOI22S $T=1001920 1071960 0 180 $X=998200 $Y=1066540
X3156 5903 5870 5902 1081 1 5865 2 AOI22S $T=1002540 940920 1 180 $X=998820 $Y=940540
X3157 5903 5870 5899 5823 1 5855 2 AOI22S $T=1003160 971160 1 180 $X=999440 $Y=970780
X3158 5883 5887 5898 5791 1 5805 2 AOI22S $T=1003160 1021560 1 180 $X=999440 $Y=1021180
X3159 5903 5870 5904 5893 1 5890 2 AOI22S $T=1003780 991320 1 180 $X=1000060 $Y=990940
X3160 5883 5887 5916 5820 1 1085 2 AOI22S $T=1003780 1041720 1 180 $X=1000060 $Y=1041340
X3161 5920 5901 1103 1094 1 5889 2 AOI22S $T=1004400 900600 1 180 $X=1000680 $Y=900220
X3162 5903 5870 5906 1079 1 5874 2 AOI22S $T=1004400 961080 0 180 $X=1000680 $Y=955660
X3163 5892 5877 5896 1095 1 1098 2 AOI22S $T=1000680 1082040 0 0 $X=1000680 $Y=1081660
X3164 5920 5901 1101 5885 1 5824 2 AOI22S $T=1005640 910680 0 180 $X=1001920 $Y=905260
X3165 5892 5877 5925 5934 1 1111 2 AOI22S $T=1004400 1071960 0 0 $X=1004400 $Y=1071580
X3166 5920 5901 1107 5819 1 1106 2 AOI22S $T=1005640 910680 0 0 $X=1005640 $Y=910300
X3167 5962 5937 5947 5960 1 5932 2 AOI22S $T=1013700 1011480 0 180 $X=1009980 $Y=1006060
X3168 1116 5937 5948 5965 1 5963 2 AOI22S $T=1009980 1051800 1 0 $X=1009980 $Y=1046380
X3169 5962 5937 5973 5929 1 5836 2 AOI22S $T=1014320 971160 1 180 $X=1010600 $Y=970780
X3170 5962 5937 5936 5974 1 5884 2 AOI22S $T=1011220 1021560 1 0 $X=1011220 $Y=1016140
X3171 5920 5968 5978 1088 1 5886 2 AOI22S $T=1015560 930840 1 180 $X=1011840 $Y=930460
X3172 5962 5968 5984 5982 1 1133 2 AOI22S $T=1014940 961080 1 0 $X=1014940 $Y=955660
X3173 1137 1134 6003 6025 1 5957 2 AOI22S $T=1018660 961080 1 0 $X=1018660 $Y=955660
X3174 6010 1134 5991 5996 1 6019 2 AOI22S $T=1018660 981240 1 0 $X=1018660 $Y=975820
X3175 6010 1140 5944 6017 1 6015 2 AOI22S $T=1022380 1041720 0 180 $X=1018660 $Y=1036300
X3176 1137 1134 6006 1141 1 1143 2 AOI22S $T=1019280 940920 0 0 $X=1019280 $Y=940540
X3177 6010 1134 5959 6023 1 1144 2 AOI22S $T=1019280 991320 1 0 $X=1019280 $Y=985900
X3178 5920 5901 1139 5987 1 6012 2 AOI22S $T=1019900 910680 0 0 $X=1019900 $Y=910300
X3179 6010 1140 5928 6032 1 6036 2 AOI22S $T=1021760 1021560 1 0 $X=1021760 $Y=1016140
X3180 6010 6004 5943 6035 1 6040 2 AOI22S $T=1022380 1011480 1 0 $X=1022380 $Y=1006060
X3181 6108 6130 5995 6009 1 6122 2 AOI22S $T=1044080 991320 0 180 $X=1040360 $Y=985900
X3182 6108 6113 5956 6138 1 6143 2 AOI22S $T=1042220 991320 0 0 $X=1042220 $Y=990940
X3183 6108 6113 5939 6132 1 1172 2 AOI22S $T=1042220 1011480 0 0 $X=1042220 $Y=1011100
X3184 1168 1165 5977 6134 1 1174 2 AOI22S $T=1043460 1061880 0 0 $X=1043460 $Y=1061500
X3185 6141 1173 6013 1171 1 6074 2 AOI22S $T=1044700 951000 1 0 $X=1044700 $Y=945580
X3186 5920 6153 1170 6135 1 6159 2 AOI22S $T=1045320 900600 0 0 $X=1045320 $Y=900220
X3187 6141 6130 6008 6149 1 1178 2 AOI22S $T=1045320 971160 1 0 $X=1045320 $Y=965740
X3188 6191 6169 6174 5990 1 6139 2 AOI22S $T=1053380 940920 1 180 $X=1049660 $Y=940540
X3189 1116 6153 6183 6165 1 1184 2 AOI22S $T=1058960 930840 1 180 $X=1055240 $Y=930460
X3190 6078 6199 6175 6171 1 6203 2 AOI22S $T=1056480 971160 1 0 $X=1056480 $Y=965740
X3191 1116 6153 6205 6213 1 1202 2 AOI22S $T=1058960 930840 0 0 $X=1058960 $Y=930460
X3192 6141 6130 6173 6210 1 6225 2 AOI22S $T=1059580 991320 1 0 $X=1059580 $Y=985900
X3193 1168 1165 1200 6228 1 1206 2 AOI22S $T=1060200 1071960 1 0 $X=1060200 $Y=1066540
X3194 1204 6153 1205 6237 1 6246 2 AOI22S $T=1062060 900600 0 0 $X=1062060 $Y=900220
X3195 6191 6169 6212 6251 1 6244 2 AOI22S $T=1062060 940920 0 0 $X=1062060 $Y=940540
X3196 6141 6130 6233 6224 1 6248 2 AOI22S $T=1062680 971160 0 0 $X=1062680 $Y=970780
X3197 6287 6199 6226 6232 1 1211 2 AOI22S $T=1073840 961080 0 180 $X=1070120 $Y=955660
X3198 6141 6130 6280 6260 1 6294 2 AOI22S $T=1071980 971160 0 0 $X=1071980 $Y=970780
X3199 6287 6199 6288 1213 1 6298 2 AOI22S $T=1074460 961080 1 0 $X=1074460 $Y=955660
X3200 6192 6277 6323 6221 1 6220 2 AOI22S $T=1080660 1051800 0 180 $X=1076940 $Y=1046380
X3201 6321 6277 1225 1215 1 6267 2 AOI22S $T=1081280 1071960 0 180 $X=1077560 $Y=1066540
X3202 6191 6169 6325 6343 1 1233 2 AOI22S $T=1084380 940920 0 0 $X=1084380 $Y=940540
X3203 6321 6338 6349 6339 1 6293 2 AOI22S $T=1088100 1071960 0 180 $X=1084380 $Y=1066540
X3204 6321 6338 6352 6322 1 6257 2 AOI22S $T=1088720 1061880 1 180 $X=1085000 $Y=1061500
X3205 6342 6348 6313 6320 1 6350 2 AOI22S $T=1086240 930840 1 0 $X=1086240 $Y=925420
X3206 6192 6169 6369 1226 1 1219 2 AOI22S $T=1089960 1001400 0 180 $X=1086240 $Y=995980
X3207 1243 6378 6389 6360 1 6311 2 AOI22S $T=1096780 1031640 0 180 $X=1093060 $Y=1026220
X3208 6342 6378 6388 6328 1 6376 2 AOI22S $T=1097400 1001400 1 180 $X=1093680 $Y=1001020
X3209 6191 6169 6390 6344 1 6381 2 AOI22S $T=1094920 951000 1 0 $X=1094920 $Y=945580
X3210 6191 6169 6391 6351 1 6371 2 AOI22S $T=1094920 971160 0 0 $X=1094920 $Y=970780
X3211 6416 6304 6380 1237 1 1231 2 AOI22S $T=1099880 1061880 1 180 $X=1096160 $Y=1061500
X3212 1256 6412 6382 6386 1 1248 2 AOI22S $T=1100500 1071960 0 180 $X=1096780 $Y=1066540
X3213 6342 6378 6409 6414 1 1255 2 AOI22S $T=1097400 981240 0 0 $X=1097400 $Y=980860
X3214 1260 1241 1259 1254 1 1253 2 AOI22S $T=1102360 910680 0 180 $X=1098640 $Y=905260
X3215 6287 6412 6397 6331 1 6427 2 AOI22S $T=1099260 1031640 0 0 $X=1099260 $Y=1031260
X3216 6287 6412 6401 6411 1 6421 2 AOI22S $T=1103600 1021560 0 180 $X=1099880 $Y=1016140
X3217 6342 6348 6424 6430 1 6413 2 AOI22S $T=1101120 930840 1 0 $X=1101120 $Y=925420
X3218 1256 6412 6425 6395 1 6436 2 AOI22S $T=1101120 1071960 1 0 $X=1101120 $Y=1066540
X3219 6416 6304 6434 6418 1 6448 2 AOI22S $T=1103600 1061880 1 0 $X=1103600 $Y=1056460
X3220 6440 1247 6419 6452 1 1262 2 AOI22S $T=1104220 971160 1 0 $X=1104220 $Y=965740
X3221 6287 6412 6396 6453 1 6405 2 AOI22S $T=1105460 1001400 1 0 $X=1105460 $Y=995980
X3222 6416 6304 6451 6446 1 6469 2 AOI22S $T=1107320 1061880 1 0 $X=1107320 $Y=1056460
X3223 1260 6348 1276 6457 1 6485 2 AOI22S $T=1109800 920760 1 0 $X=1109800 $Y=915340
X3224 6416 1173 6402 6501 1 6506 2 AOI22S $T=1114140 991320 0 0 $X=1114140 $Y=990940
X3225 6223 1173 6422 6513 1 6500 2 AOI22S $T=1119720 971160 0 0 $X=1119720 $Y=970780
X3226 3745 3751 3756 3761 2 1 3777 AN4S $T=625580 981240 1 0 $X=625580 $Y=975820
X3227 3781 3783 3788 3773 2 1 3803 AN4S $T=631780 981240 1 0 $X=631780 $Y=975820
X3228 3802 3796 3799 3814 2 1 3826 AN4S $T=637980 981240 1 0 $X=637980 $Y=975820
X3229 3892 3879 3932 3910 2 1 3966 AN4S $T=661540 961080 0 0 $X=661540 $Y=960700
X3230 3928 3930 3913 3882 2 1 3955 AN4S $T=661540 971160 1 0 $X=661540 $Y=965740
X3231 4044 4038 4031 4028 2 1 4018 AN4S $T=680140 971160 0 180 $X=675180 $Y=965740
X3232 4083 4082 4059 4070 2 1 4032 AN4S $T=686960 961080 1 180 $X=682000 $Y=960700
X3233 4145 4138 3868 4067 2 1 646 AN4S $T=697500 920760 0 180 $X=692540 $Y=915340
X3234 4174 4168 3921 4074 2 1 649 AN4S $T=701840 910680 0 180 $X=696880 $Y=905260
X3235 4242 4243 4237 4234 2 1 4175 AN4S $T=714860 961080 0 180 $X=709900 $Y=955660
X3236 4292 4286 4274 4249 2 1 4256 AN4S $T=724160 971160 1 180 $X=719200 $Y=970780
X3237 4330 4327 4302 4222 2 1 4296 AN4S $T=729120 971160 0 180 $X=724160 $Y=965740
X3238 5278 926 5266 5110 2 1 920 AN4S $T=886600 900600 1 180 $X=881640 $Y=900220
X3239 5279 5240 5267 5014 2 1 921 AN4S $T=886600 910680 1 180 $X=881640 $Y=910300
X3240 5257 5254 5271 5066 2 1 931 AN4S $T=882880 920760 1 0 $X=882880 $Y=915340
X3241 5292 5251 5303 5120 2 1 936 AN4S $T=887220 910680 0 0 $X=887220 $Y=910300
X3242 5898 5936 5928 5923 2 1 5620 AN4S $T=1008120 1021560 1 180 $X=1003160 $Y=1021180
X3243 5879 5947 5943 5939 2 1 5614 AN4S $T=1009980 1011480 0 180 $X=1005020 $Y=1006060
X3244 5916 5948 5944 5940 2 1 5586 AN4S $T=1009980 1041720 1 180 $X=1005020 $Y=1041340
X3245 5896 1114 1112 5942 2 1 5495 AN4S $T=1009980 1082040 1 180 $X=1005020 $Y=1081660
X3246 5904 5969 5959 5956 2 1 5632 AN4S $T=1013700 1001400 0 180 $X=1008740 $Y=995980
X3247 5891 5952 5971 5977 2 1 5477 AN4S $T=1010600 1061880 0 0 $X=1010600 $Y=1061500
X3248 5899 5973 5991 5995 2 1 5552 AN4S $T=1014320 971160 0 0 $X=1014320 $Y=970780
X3249 5906 5984 6003 6008 2 1 5601 AN4S $T=1016180 951000 0 0 $X=1016180 $Y=950620
X3250 5902 5978 6006 6013 2 1 5519 AN4S $T=1016800 951000 1 0 $X=1016800 $Y=945580
X3251 6174 6183 6175 6173 2 1 5708 AN4S $T=1055240 971160 0 180 $X=1050280 $Y=965740
X3252 6212 6205 6226 6233 2 1 5625 AN4S $T=1060820 961080 1 0 $X=1060820 $Y=955660
X3253 6325 6313 6288 6280 2 1 5787 AN4S $T=1081900 951000 1 180 $X=1076940 $Y=950620
X3254 6349 1246 6382 6380 2 1 5714 AN4S $T=1096780 1071960 0 180 $X=1091820 $Y=1066540
X3255 6369 6388 6396 6402 2 1 5752 AN4S $T=1094300 1001400 1 0 $X=1094300 $Y=995980
X3256 6292 6389 6397 6403 2 1 5690 AN4S $T=1094300 1031640 0 0 $X=1094300 $Y=1031260
X3257 6305 6379 6401 6407 2 1 5720 AN4S $T=1094920 1021560 1 0 $X=1094920 $Y=1016140
X3258 6391 6409 6419 6422 2 1 5735 AN4S $T=1098640 971160 1 0 $X=1098640 $Y=965740
X3259 6323 1257 6425 6434 2 1 5745 AN4S $T=1099880 1051800 1 0 $X=1099880 $Y=1046380
X3260 6390 6424 6431 6435 2 1 5762 AN4S $T=1101120 951000 1 0 $X=1101120 $Y=945580
X3261 6352 1272 6454 6451 2 1 5713 AN4S $T=1109800 1061880 1 180 $X=1104840 $Y=1061500
X3262 33 2 1 1550 BUF1 $T=254820 900600 0 0 $X=254820 $Y=900220
X3263 1820 2 1 1538 BUF1 $T=297600 1031640 0 180 $X=295120 $Y=1026220
X3264 69 2 1 1790 BUF1 $T=302560 930840 0 0 $X=302560 $Y=930460
X3265 99 2 1 1880 BUF1 $T=313720 951000 1 180 $X=311240 $Y=950620
X3266 96 2 1 1868 BUF1 $T=326740 920760 0 0 $X=326740 $Y=920380
X3267 139 2 1 2071 BUF1 $T=337900 930840 0 0 $X=337900 $Y=930460
X3268 198 2 1 2402 BUF1 $T=382540 1082040 1 0 $X=382540 $Y=1076620
X3269 2483 2 1 208 BUF1 $T=399900 1071960 1 180 $X=397420 $Y=1071580
X3270 2419 2 1 2523 BUF1 $T=404240 1041720 0 0 $X=404240 $Y=1041340
X3271 2539 2 1 2433 BUF1 $T=411680 1041720 1 180 $X=409200 $Y=1041340
X3272 2624 2 1 2535 BUF1 $T=420360 1071960 1 180 $X=417880 $Y=1071580
X3273 2624 2 1 239 BUF1 $T=422220 1082040 1 180 $X=419740 $Y=1081660
X3274 2539 2 1 2680 BUF1 $T=429040 1031640 0 0 $X=429040 $Y=1031260
X3275 249 2 1 2702 BUF1 $T=430280 900600 0 0 $X=430280 $Y=900220
X3276 2483 2 1 254 BUF1 $T=432140 1071960 0 0 $X=432140 $Y=1071580
X3277 2721 2 1 2556 BUF1 $T=443300 1041720 1 0 $X=443300 $Y=1036300
X3278 2624 2 1 2793 BUF1 $T=451360 1031640 0 0 $X=451360 $Y=1031260
X3279 2454 2 1 284 BUF1 $T=453220 1071960 0 0 $X=453220 $Y=1071580
X3280 285 2 1 198 BUF1 $T=461280 1082040 1 180 $X=458800 $Y=1081660
X3281 297 2 1 2650 BUF1 $T=466240 940920 1 180 $X=463760 $Y=940540
X3282 295 2 1 2747 BUF1 $T=466240 951000 0 180 $X=463760 $Y=945580
X3283 2884 2 1 2768 BUF1 $T=467480 971160 1 180 $X=465000 $Y=970780
X3284 277 2 1 2888 BUF1 $T=465620 920760 0 0 $X=465620 $Y=920380
X3285 2908 2 1 2579 BUF1 $T=476160 981240 0 0 $X=476160 $Y=980860
X3286 311 2 1 2721 BUF1 $T=484220 991320 0 180 $X=481740 $Y=985900
X3287 2997 2 1 2818 BUF1 $T=484220 1031640 0 180 $X=481740 $Y=1026220
X3288 314 2 1 2624 BUF1 $T=485460 981240 0 180 $X=482980 $Y=975820
X3289 2990 2 1 2819 BUF1 $T=486700 1051800 1 180 $X=484220 $Y=1051420
X3290 3004 2 1 306 BUF1 $T=491040 1071960 1 0 $X=491040 $Y=1066540
X3291 2702 2 1 3053 BUF1 $T=494140 920760 0 0 $X=494140 $Y=920380
X3292 3059 2 1 310 BUF1 $T=497860 1071960 0 0 $X=497860 $Y=1071580
X3293 3067 2 1 2992 BUF1 $T=502820 951000 0 180 $X=500340 $Y=945580
X3294 332 2 1 3059 BUF1 $T=502820 1011480 0 0 $X=502820 $Y=1011100
X3295 343 2 1 289 BUF1 $T=507160 910680 1 180 $X=504680 $Y=910300
X3296 340 2 1 2483 BUF1 $T=507160 930840 1 180 $X=504680 $Y=930460
X3297 331 2 1 351 BUF1 $T=510880 910680 0 0 $X=510880 $Y=910300
X3298 352 2 1 3123 BUF1 $T=514600 910680 0 180 $X=512120 $Y=905260
X3299 295 2 1 3175 BUF1 $T=519560 940920 0 0 $X=519560 $Y=940540
X3300 3176 2 1 2997 BUF1 $T=522040 1031640 0 180 $X=519560 $Y=1026220
X3301 3192 2 1 3177 BUF1 $T=522660 1051800 0 0 $X=522660 $Y=1051420
X3302 363 2 1 2906 BUF1 $T=526380 951000 0 180 $X=523900 $Y=945580
X3303 3079 2 1 3115 BUF1 $T=524520 1031640 1 0 $X=524520 $Y=1026220
X3304 3233 2 1 3166 BUF1 $T=530720 971160 1 180 $X=528240 $Y=970780
X3305 183 2 1 3079 BUF1 $T=528240 1041720 1 0 $X=528240 $Y=1036300
X3306 297 2 1 3280 BUF1 $T=536920 940920 0 0 $X=536920 $Y=940540
X3307 363 2 1 3113 BUF1 $T=536920 951000 0 0 $X=536920 $Y=950620
X3308 2888 2 1 3276 BUF1 $T=536920 1051800 0 0 $X=536920 $Y=1051420
X3309 3271 2 1 3185 BUF1 $T=537540 1051800 1 0 $X=537540 $Y=1046380
X3310 3079 2 1 3306 BUF1 $T=541880 1031640 0 0 $X=541880 $Y=1031260
X3311 403 2 1 3233 BUF1 $T=547460 940920 1 180 $X=544980 $Y=940540
X3312 388 2 1 3176 BUF1 $T=553660 910680 0 180 $X=551180 $Y=905260
X3313 3203 2 1 415 BUF1 $T=551180 940920 0 0 $X=551180 $Y=940540
X3314 3359 2 1 3217 BUF1 $T=557380 971160 0 180 $X=554900 $Y=965740
X3315 2902 2 1 3401 BUF1 $T=558620 920760 0 0 $X=558620 $Y=920380
X3316 3175 2 1 3420 BUF1 $T=571020 961080 0 180 $X=568540 $Y=955660
X3317 407 2 1 3443 BUF1 $T=572880 971160 1 0 $X=572880 $Y=965740
X3318 294 2 1 3492 BUF1 $T=575980 910680 0 0 $X=575980 $Y=910300
X3319 2790 2 1 460 BUF1 $T=579080 1082040 1 0 $X=579080 $Y=1076620
X3320 3271 2 1 3396 BUF1 $T=580320 1061880 1 0 $X=580320 $Y=1056460
X3321 3500 2 1 3400 BUF1 $T=583420 1021560 1 0 $X=583420 $Y=1016140
X3322 473 2 1 3271 BUF1 $T=585900 1001400 1 0 $X=585900 $Y=995980
X3323 451 2 1 3500 BUF1 $T=590240 940920 1 180 $X=587760 $Y=940540
X3324 3053 2 1 3556 BUF1 $T=590240 920760 1 0 $X=590240 $Y=915340
X3325 407 2 1 484 BUF1 $T=594580 920760 0 0 $X=594580 $Y=920380
X3326 3654 2 1 3359 BUF1 $T=615660 971160 0 180 $X=613180 $Y=965740
X3327 3401 2 1 3722 BUF1 $T=618760 920760 0 0 $X=618760 $Y=920380
X3328 3620 2 1 3687 BUF1 $T=624340 1031640 1 180 $X=621860 $Y=1031260
X3329 3556 2 1 3747 BUF1 $T=636120 920760 1 180 $X=633640 $Y=920380
X3330 3276 2 1 543 BUF1 $T=635500 1061880 1 0 $X=635500 $Y=1056460
X3331 3836 2 1 3674 BUF1 $T=646040 1061880 0 180 $X=643560 $Y=1056460
X3332 3280 2 1 3846 BUF1 $T=644800 961080 1 0 $X=644800 $Y=955660
X3333 3832 2 1 3656 BUF1 $T=648520 1061880 0 180 $X=646040 $Y=1056460
X3334 3556 2 1 3854 BUF1 $T=646660 920760 1 0 $X=646660 $Y=915340
X3335 585 2 1 572 BUF1 $T=663400 900600 1 180 $X=660920 $Y=900220
X3336 534 2 1 598 BUF1 $T=666500 1082040 0 0 $X=666500 $Y=1081660
X3337 3316 2 1 588 BUF1 $T=669600 940920 1 180 $X=667120 $Y=940540
X3338 3587 2 1 3987 BUF1 $T=673320 1021560 1 0 $X=673320 $Y=1016140
X3339 598 2 1 627 BUF1 $T=678900 1082040 0 0 $X=678900 $Y=1081660
X3340 3987 2 1 3969 BUF1 $T=680140 1041720 0 0 $X=680140 $Y=1041340
X3341 3891 2 1 643 BUF1 $T=685720 1082040 1 0 $X=685720 $Y=1076620
X3342 3697 2 1 4103 BUF1 $T=686340 1041720 1 0 $X=686340 $Y=1036300
X3343 3722 2 1 4132 BUF1 $T=693160 910680 1 0 $X=693160 $Y=905260
X3344 4139 2 1 3836 BUF1 $T=697500 1051800 0 180 $X=695020 $Y=1046380
X3345 663 2 1 4226 BUF1 $T=709280 920760 0 0 $X=709280 $Y=920380
X3346 4226 2 1 4008 BUF1 $T=712380 991320 0 180 $X=709900 $Y=985900
X3347 3846 2 1 4250 BUF1 $T=719200 1001400 1 0 $X=719200 $Y=995980
X3348 4310 2 1 4078 BUF1 $T=725400 1001400 1 180 $X=722920 $Y=1001020
X3349 4139 2 1 4315 BUF1 $T=724160 1051800 0 0 $X=724160 $Y=1051420
X3350 4310 2 1 4139 BUF1 $T=725400 1001400 1 0 $X=725400 $Y=995980
X3351 4158 2 1 4100 BUF1 $T=726020 1011480 1 0 $X=726020 $Y=1006060
X3352 4328 2 1 4158 BUF1 $T=729120 991320 1 180 $X=726640 $Y=990940
X3353 694 2 1 4328 BUF1 $T=733460 910680 0 180 $X=730980 $Y=905260
X3354 702 2 1 4310 BUF1 $T=735940 910680 0 180 $X=733460 $Y=905260
X3355 3834 2 1 4380 BUF1 $T=737800 971160 1 0 $X=737800 $Y=965740
X3356 705 2 1 711 BUF1 $T=741520 1051800 0 0 $X=741520 $Y=1051420
X3357 4380 2 1 4421 BUF1 $T=746480 1011480 1 0 $X=746480 $Y=1006060
X3358 4340 2 1 4444 BUF1 $T=748340 1031640 0 0 $X=748340 $Y=1031260
X3359 721 2 1 4454 BUF1 $T=750200 920760 0 0 $X=750200 $Y=920380
X3360 722 2 1 3994 BUF1 $T=750200 940920 0 0 $X=750200 $Y=940540
X3361 709 2 1 4413 BUF1 $T=752680 1061880 1 180 $X=750200 $Y=1061500
X3362 4441 2 1 4533 BUF1 $T=766320 961080 1 0 $X=766320 $Y=955660
X3363 4533 2 1 4542 BUF1 $T=766320 1041720 0 0 $X=766320 $Y=1041340
X3364 4250 2 1 4520 BUF1 $T=766940 1011480 0 0 $X=766940 $Y=1011100
X3365 4576 2 1 4555 BUF1 $T=774380 971160 1 180 $X=771900 $Y=970780
X3366 4378 2 1 4609 BUF1 $T=773140 981240 1 0 $X=773140 $Y=975820
X3367 752 2 1 4146 BUF1 $T=773760 920760 0 0 $X=773760 $Y=920380
X3368 4597 2 1 4540 BUF1 $T=776860 951000 1 180 $X=774380 $Y=950620
X3369 4600 2 1 4576 BUF1 $T=777480 940920 1 180 $X=775000 $Y=940540
X3370 4557 2 1 754 BUF1 $T=778720 1061880 1 180 $X=776240 $Y=1061500
X3371 4132 2 1 4623 BUF1 $T=776860 981240 0 0 $X=776860 $Y=980860
X3372 763 2 1 4579 BUF1 $T=778100 900600 0 0 $X=778100 $Y=900220
X3373 723 2 1 4635 BUF1 $T=779340 930840 0 0 $X=779340 $Y=930460
X3374 782 2 1 709 BUF1 $T=786160 1082040 0 180 $X=783680 $Y=1076620
X3375 4727 2 1 796 BUF1 $T=796080 1082040 0 180 $X=793600 $Y=1076620
X3376 4782 2 1 4686 BUF1 $T=804140 981240 1 180 $X=801660 $Y=980860
X3377 4823 2 1 4782 BUF1 $T=812820 951000 1 180 $X=810340 $Y=950620
X3378 4848 2 1 822 BUF1 $T=811580 1071960 0 0 $X=811580 $Y=1071580
X3379 779 2 1 4727 BUF1 $T=813440 1071960 1 0 $X=813440 $Y=1066540
X3380 4861 2 1 835 BUF1 $T=814060 900600 0 0 $X=814060 $Y=900220
X3381 832 2 1 4813 BUF1 $T=816540 951000 1 180 $X=814060 $Y=950620
X3382 782 2 1 841 BUF1 $T=817160 1082040 1 0 $X=817160 $Y=1076620
X3383 4542 2 1 4911 BUF1 $T=820880 1041720 1 0 $X=820880 $Y=1036300
X3384 832 2 1 4924 BUF1 $T=823980 951000 1 0 $X=823980 $Y=945580
X3385 4131 2 1 4934 BUF1 $T=826460 1061880 1 0 $X=826460 $Y=1056460
X3386 4883 2 1 823 BUF1 $T=829560 1041720 0 180 $X=827080 $Y=1036300
X3387 856 2 1 4823 BUF1 $T=830800 920760 1 180 $X=828320 $Y=920380
X3388 4520 2 1 4968 BUF1 $T=832660 1031640 1 0 $X=832660 $Y=1026220
X3389 863 2 1 4597 BUF1 $T=835140 920760 0 0 $X=835140 $Y=920380
X3390 4444 2 1 4982 BUF1 $T=835140 1041720 0 0 $X=835140 $Y=1041340
X3391 4600 2 1 4997 BUF1 $T=837620 951000 1 0 $X=837620 $Y=945580
X3392 4597 2 1 4992 BUF1 $T=843200 951000 1 180 $X=840720 $Y=950620
X3393 4848 2 1 883 BUF1 $T=851260 1071960 1 0 $X=851260 $Y=1066540
X3394 5086 2 1 5034 BUF1 $T=856840 961080 1 180 $X=854360 $Y=960700
X3395 5055 2 1 886 BUF1 $T=854360 1061880 0 0 $X=854360 $Y=1061500
X3396 5081 2 1 5086 BUF1 $T=854980 971160 1 0 $X=854980 $Y=965740
X3397 4623 2 1 5081 BUF1 $T=857460 981240 1 180 $X=854980 $Y=980860
X3398 4454 2 1 5070 BUF1 $T=859320 1001400 1 0 $X=859320 $Y=995980
X3399 4727 2 1 901 BUF1 $T=864280 1061880 0 0 $X=864280 $Y=1061500
X3400 4635 2 1 5262 BUF1 $T=881640 971160 0 0 $X=881640 $Y=970780
X3401 4533 2 1 5258 BUF1 $T=883500 961080 1 0 $X=883500 $Y=955660
X3402 4579 2 1 5264 BUF1 $T=883500 1031640 0 0 $X=883500 $Y=1031260
X3403 5214 2 1 925 BUF1 $T=886600 1071960 1 0 $X=886600 $Y=1066540
X3404 5050 2 1 5315 BUF1 $T=887220 991320 1 0 $X=887220 $Y=985900
X3405 5264 2 1 923 BUF1 $T=890320 1061880 1 180 $X=887840 $Y=1061500
X3406 5086 2 1 948 BUF1 $T=897760 910680 0 0 $X=897760 $Y=910300
X3407 4623 2 1 5395 BUF1 $T=902720 1041720 1 0 $X=902720 $Y=1036300
X3408 969 2 1 5433 BUF1 $T=913260 1082040 1 0 $X=913260 $Y=1076620
X3409 485 2 1 987 BUF1 $T=920700 920760 0 0 $X=920700 $Y=920380
X3410 5258 2 1 5500 BUF1 $T=924420 1011480 1 0 $X=924420 $Y=1006060
X3411 4854 2 1 5486 BUF1 $T=927520 961080 0 0 $X=927520 $Y=960700
X3412 1000 2 1 5534 BUF1 $T=930000 900600 0 0 $X=930000 $Y=900220
X3413 1007 2 1 5526 BUF1 $T=934340 961080 1 0 $X=934340 $Y=955660
X3414 5545 2 1 5465 BUF1 $T=934960 1041720 0 0 $X=934960 $Y=1041340
X3415 1012 2 1 5496 BUF1 $T=939300 961080 0 180 $X=936820 $Y=955660
X3416 1012 2 1 5594 BUF1 $T=940540 940920 1 0 $X=940540 $Y=935500
X3417 5534 2 1 1028 BUF1 $T=950460 961080 1 0 $X=950460 $Y=955660
X3418 5465 2 1 5655 BUF1 $T=952320 1061880 0 0 $X=952320 $Y=1061500
X3419 5559 2 1 5644 BUF1 $T=961620 1041720 1 0 $X=961620 $Y=1036300
X3420 5258 2 1 5729 BUF1 $T=962860 971160 0 0 $X=962860 $Y=970780
X3421 1052 2 1 5559 BUF1 $T=965960 1011480 1 180 $X=963480 $Y=1011100
X3422 5395 2 1 1059 BUF1 $T=964100 1071960 0 0 $X=964100 $Y=1071580
X3423 5262 2 1 5821 BUF1 $T=981460 1051800 0 0 $X=981460 $Y=1051420
X3424 5821 2 1 5777 BUF1 $T=985800 1051800 0 0 $X=985800 $Y=1051420
X3425 1090 2 1 5866 BUF1 $T=998820 930840 0 0 $X=998820 $Y=930460
X3426 1091 2 1 5883 BUF1 $T=998820 940920 1 0 $X=998820 $Y=935500
X3427 5887 2 1 5877 BUF1 $T=1000680 1071960 0 0 $X=1000680 $Y=1071580
X3428 5883 2 1 5892 BUF1 $T=1002540 1071960 1 0 $X=1002540 $Y=1066540
X3429 5937 2 1 1113 BUF1 $T=1006260 1051800 1 0 $X=1006260 $Y=1046380
X3430 929 2 1 1099 BUF1 $T=1006880 971160 0 0 $X=1006880 $Y=970780
X3431 5968 2 1 5937 BUF1 $T=1013700 961080 0 180 $X=1011220 $Y=955660
X3432 1125 2 1 1116 BUF1 $T=1014320 930840 0 180 $X=1011840 $Y=925420
X3433 6010 2 1 1148 BUF1 $T=1023620 1051800 0 0 $X=1023620 $Y=1051420
X3434 5486 2 1 6039 BUF1 $T=1024240 951000 1 0 $X=1024240 $Y=945580
X3435 1162 2 1 5968 BUF1 $T=1037880 910680 1 0 $X=1037880 $Y=905260
X3436 5821 2 1 5976 BUF1 $T=1039120 1051800 1 0 $X=1039120 $Y=1046380
X3437 6108 2 1 1168 BUF1 $T=1040980 1061880 0 0 $X=1040980 $Y=1061500
X3438 6141 2 1 6108 BUF1 $T=1047180 991320 0 180 $X=1044700 $Y=985900
X3439 6130 2 1 6113 BUF1 $T=1045940 991320 0 0 $X=1045940 $Y=990940
X3440 841 2 1 1182 BUF1 $T=1046560 1082040 1 0 $X=1046560 $Y=1076620
X3441 6113 2 1 1165 BUF1 $T=1047180 1061880 0 0 $X=1047180 $Y=1061500
X3442 1091 2 1 6192 BUF1 $T=1053380 940920 0 0 $X=1053380 $Y=940540
X3443 6101 2 1 6206 BUF1 $T=1062680 961080 0 0 $X=1062680 $Y=960700
X3444 6071 2 1 6315 BUF1 $T=1080040 930840 1 0 $X=1080040 $Y=925420
X3445 1176 2 1 6330 BUF1 $T=1080040 1021560 1 0 $X=1080040 $Y=1016140
X3446 6315 2 1 6299 BUF1 $T=1083140 951000 0 180 $X=1080660 $Y=945580
X3447 1125 2 1 6342 BUF1 $T=1082520 920760 1 0 $X=1082520 $Y=915340
X3448 1162 2 1 6348 BUF1 $T=1084380 910680 0 0 $X=1084380 $Y=910300
X3449 6097 2 1 1239 BUF1 $T=1088100 1071960 1 0 $X=1088100 $Y=1066540
X3450 1221 2 1 1238 BUF1 $T=1088720 1061880 0 0 $X=1088720 $Y=1061500
X3451 6342 2 1 1243 BUF1 $T=1095540 1011480 1 180 $X=1093060 $Y=1011100
X3452 1252 2 1 6378 BUF1 $T=1100500 1021560 1 180 $X=1098020 $Y=1021180
X3453 6342 2 1 1260 BUF1 $T=1101740 920760 1 0 $X=1101740 $Y=915340
X3454 1256 2 1 6287 BUF1 $T=1102360 1001400 1 0 $X=1102360 $Y=995980
X3455 6060 2 1 6426 BUF1 $T=1105460 981240 1 0 $X=1105460 $Y=975820
X3456 6348 2 1 1252 BUF1 $T=1108560 930840 0 180 $X=1106080 $Y=925420
X3457 1274 2 1 1273 BUF1 $T=1111040 930840 1 180 $X=1108560 $Y=930460
X3458 5821 2 1 1266 BUF1 $T=1111660 1071960 0 180 $X=1109180 $Y=1066540
X3459 6223 2 1 6416 BUF1 $T=1115380 971160 0 0 $X=1115380 $Y=970780
X3460 1265 2 1 6366 BUF1 $T=1122820 930840 0 0 $X=1122820 $Y=930460
X3461 48 1 2 61 BUF1CK $T=274040 900600 0 0 $X=274040 $Y=900220
X3462 1657 1 2 1826 BUF1CK $T=295120 1011480 0 0 $X=295120 $Y=1011100
X3463 83 1 2 1895 BUF1CK $T=304420 991320 1 0 $X=304420 $Y=985900
X3464 92 1 2 1922 BUF1CK $T=309380 1001400 0 0 $X=309380 $Y=1001020
X3465 1923 1 2 1929 BUF1CK $T=310620 1021560 1 0 $X=310620 $Y=1016140
X3466 1807 1 2 1865 BUF1CK $T=314340 1001400 0 0 $X=314340 $Y=1001020
X3467 123 1 2 2011 BUF1CK $T=324880 1021560 0 0 $X=324880 $Y=1021180
X3468 2097 1 2 2108 BUF1CK $T=337900 1061880 1 0 $X=337900 $Y=1056460
X3469 1849 1 2 2097 BUF1CK $T=342240 1051800 0 0 $X=342240 $Y=1051420
X3470 2556 1 2 2419 BUF1CK $T=411060 1051800 0 180 $X=408580 $Y=1046380
X3471 2600 1 2 2605 BUF1CK $T=416020 961080 1 0 $X=416020 $Y=955660
X3472 2676 1 2 2652 BUF1CK $T=432760 1031640 1 0 $X=432760 $Y=1026220
X3473 2728 1 2 211 BUF1CK $T=441440 1082040 0 180 $X=438960 $Y=1076620
X3474 2892 1 2 2903 BUF1CK $T=468100 1001400 1 0 $X=468100 $Y=995980
X3475 2483 1 2 2904 BUF1CK $T=468100 1031640 0 0 $X=468100 $Y=1031260
X3476 2992 1 2 3062 BUF1CK $T=502200 971160 0 180 $X=499720 $Y=965740
X3477 3077 1 2 3004 BUF1CK $T=505300 1041720 0 180 $X=502820 $Y=1036300
X3478 3359 1 2 3067 BUF1CK $T=554900 951000 1 0 $X=554900 $Y=945580
X3479 3330 1 2 3333 BUF1CK $T=562340 951000 1 0 $X=562340 $Y=945580
X3480 3841 1 2 3696 BUF1CK $T=647900 1031640 0 180 $X=645420 $Y=1026220
X3481 3917 1 2 3926 BUF1CK $T=659060 961080 0 0 $X=659060 $Y=960700
X3482 3895 1 2 3942 BUF1CK $T=661540 951000 0 0 $X=661540 $Y=950620
X3483 4036 1 2 4045 BUF1CK $T=677660 1001400 0 0 $X=677660 $Y=1001020
X3484 4117 1 2 4122 BUF1CK $T=690680 1041720 1 0 $X=690680 $Y=1036300
X3485 4176 1 2 4183 BUF1CK $T=700600 961080 1 0 $X=700600 $Y=955660
X3486 4161 1 2 4206 BUF1CK $T=704320 1021560 0 0 $X=704320 $Y=1021180
X3487 4123 1 2 4111 BUF1CK $T=706180 1001400 1 0 $X=706180 $Y=995980
X3488 4216 1 2 4199 BUF1CK $T=711140 961080 0 0 $X=711140 $Y=960700
X3489 4259 1 2 4265 BUF1CK $T=716720 1001400 1 0 $X=716720 $Y=995980
X3490 4312 1 2 4325 BUF1CK $T=725400 961080 1 0 $X=725400 $Y=955660
X3491 4382 1 2 4384 BUF1CK $T=735320 1031640 1 0 $X=735320 $Y=1026220
X3492 4403 1 2 4400 BUF1CK $T=739660 961080 0 0 $X=739660 $Y=960700
X3493 4402 1 2 4404 BUF1CK $T=745240 920760 1 0 $X=745240 $Y=915340
X3494 4434 1 2 4445 BUF1CK $T=747720 930840 0 0 $X=747720 $Y=930460
X3495 4423 1 2 4415 BUF1CK $T=748960 1011480 1 0 $X=748960 $Y=1006060
X3496 4452 1 2 4458 BUF1CK $T=750820 930840 1 0 $X=750820 $Y=925420
X3497 4455 1 2 4464 BUF1CK $T=751440 961080 0 0 $X=751440 $Y=960700
X3498 4485 1 2 4489 BUF1CK $T=757020 1041720 1 0 $X=757020 $Y=1036300
X3499 4493 1 2 4500 BUF1CK $T=758880 1041720 0 0 $X=758880 $Y=1041340
X3500 4497 1 2 4491 BUF1CK $T=766940 930840 0 0 $X=766940 $Y=930460
X3501 4577 1 2 4588 BUF1CK $T=772520 951000 1 0 $X=772520 $Y=945580
X3502 4592 1 2 4566 BUF1CK $T=774380 981240 0 0 $X=774380 $Y=980860
X3503 4622 1 2 4618 BUF1CK $T=786160 991320 0 0 $X=786160 $Y=990940
X3504 4560 1 2 4569 BUF1CK $T=786780 920760 1 0 $X=786780 $Y=915340
X3505 4636 1 2 4556 BUF1CK $T=788020 1051800 0 0 $X=788020 $Y=1051420
X3506 4668 1 2 4667 BUF1CK $T=790500 1001400 1 0 $X=790500 $Y=995980
X3507 4763 1 2 4771 BUF1CK $T=799180 1051800 1 0 $X=799180 $Y=1046380
X3508 4757 1 2 828 BUF1CK $T=811580 900600 0 0 $X=811580 $Y=900220
X3509 825 1 2 830 BUF1CK $T=811580 910680 0 0 $X=811580 $Y=910300
X3510 4881 1 2 4892 BUF1CK $T=816540 1071960 1 0 $X=816540 $Y=1066540
X3511 789 1 2 4894 BUF1CK $T=817780 1011480 0 0 $X=817780 $Y=1011100
X3512 4742 1 2 4865 BUF1CK $T=820260 991320 0 0 $X=820260 $Y=990940
X3513 857 1 2 859 BUF1CK $T=828940 910680 1 0 $X=828940 $Y=905260
X3514 4971 1 2 4954 BUF1CK $T=835760 940920 1 0 $X=835760 $Y=935500
X3515 4910 1 2 4957 BUF1CK $T=842580 1001400 0 0 $X=842580 $Y=1001020
X3516 4944 1 2 4932 BUF1CK $T=842580 1011480 1 0 $X=842580 $Y=1006060
X3517 5085 1 2 5092 BUF1CK $T=854360 910680 0 0 $X=854360 $Y=910300
X3518 4531 1 2 5173 BUF1CK $T=867380 1021560 0 0 $X=867380 $Y=1021180
X3519 5179 1 2 5084 BUF1CK $T=875440 920760 1 0 $X=875440 $Y=915340
X3520 5079 1 2 5115 BUF1CK $T=879780 1021560 1 0 $X=879780 $Y=1016140
X3521 5313 1 2 5307 BUF1CK $T=889700 1051800 1 0 $X=889700 $Y=1046380
X3522 5352 1 2 5323 BUF1CK $T=897140 991320 1 0 $X=897140 $Y=985900
X3523 5306 1 2 5314 BUF1CK $T=899620 1061880 0 0 $X=899620 $Y=1061500
X3524 5450 1 2 5458 BUF1CK $T=919460 961080 1 0 $X=919460 $Y=955660
X3525 4966 1 2 5497 BUF1CK $T=925040 991320 0 0 $X=925040 $Y=990940
X3526 5550 1 2 5565 BUF1CK $T=935580 991320 1 0 $X=935580 $Y=985900
X3527 5643 1 2 5622 BUF1CK $T=956660 1031640 0 0 $X=956660 $Y=1031260
X3528 5650 1 2 5595 BUF1CK $T=957280 1011480 1 0 $X=957280 $Y=1006060
X3529 5696 1 2 5688 BUF1CK $T=964100 991320 0 0 $X=964100 $Y=990940
X3530 5704 1 2 5671 BUF1CK $T=969060 920760 0 0 $X=969060 $Y=920380
X3531 5839 1 2 5846 BUF1CK $T=990760 961080 0 0 $X=990760 $Y=960700
X3532 5851 1 2 5861 BUF1CK $T=992620 940920 1 0 $X=992620 $Y=935500
X3533 1120 1 2 1123 BUF1CK $T=1010600 910680 1 0 $X=1010600 $Y=905260
X3534 5961 1 2 5972 BUF1CK $T=1010600 920760 1 0 $X=1010600 $Y=915340
X3535 1128 1 2 5994 BUF1CK $T=1013700 910680 0 0 $X=1013700 $Y=910300
X3536 6028 1 2 1145 BUF1CK $T=1022380 910680 1 0 $X=1022380 $Y=905260
X3537 6007 1 2 6044 BUF1CK $T=1024860 940920 1 0 $X=1024860 $Y=935500
X3538 5809 1 2 6097 BUF1CK $T=1034160 1061880 0 0 $X=1034160 $Y=1061500
X3539 6092 1 2 6109 BUF1CK $T=1036020 1031640 1 0 $X=1036020 $Y=1026220
X3540 6148 1 2 6157 BUF1CK $T=1045320 961080 1 0 $X=1045320 $Y=955660
X3541 6096 1 2 6110 BUF1CK $T=1047180 910680 0 0 $X=1047180 $Y=910300
X3542 6083 1 2 6137 BUF1CK $T=1058340 1041720 0 0 $X=1058340 $Y=1041340
X3543 6271 1 2 6274 BUF1CK $T=1068880 910680 1 0 $X=1068880 $Y=905260
X3544 6295 1 2 6285 BUF1CK $T=1081280 910680 0 0 $X=1081280 $Y=910300
X3545 6400 1 2 6406 BUF1CK $T=1095540 1011480 0 0 $X=1095540 $Y=1011100
X3546 6227 1 2 6442 BUF1CK $T=1102980 1031640 0 0 $X=1102980 $Y=1031260
X3547 6472 1 2 6480 BUF1CK $T=1109800 1031640 1 0 $X=1109800 $Y=1026220
X3548 6492 1 2 6490 BUF1CK $T=1113520 991320 1 0 $X=1113520 $Y=985900
X3549 153 1749 1 2 INV2 $T=341620 1031640 1 180 $X=339760 $Y=1031260
X3550 434 387 1 2 INV2 $T=567300 1082040 1 180 $X=565440 $Y=1081660
X3551 3535 501 1 2 INV2 $T=605740 1051800 0 0 $X=605740 $Y=1051420
X3552 3941 3706 1 2 INV2 $T=663400 1041720 0 180 $X=661540 $Y=1036300
X3553 629 4041 1 2 INV2 $T=682620 961080 0 180 $X=680760 $Y=955660
X3554 4154 3841 1 2 INV2 $T=699360 1031640 0 180 $X=697500 $Y=1026220
X3555 662 4116 1 2 INV2 $T=726640 981240 0 0 $X=726640 $Y=980860
X3556 4134 621 1 2 INV2 $T=748340 991320 0 0 $X=748340 $Y=990940
X3557 4575 753 1 2 INV2 $T=773760 1082040 1 0 $X=773760 $Y=1076620
X3558 4075 4703 1 2 INV2 $T=792360 910680 1 0 $X=792360 $Y=905260
X3559 4830 4883 1 2 INV2 $T=821500 920760 1 0 $X=821500 $Y=915340
X3560 5656 1031 1 2 INV2 $T=954800 991320 0 0 $X=954800 $Y=990940
X3561 6002 1140 1 2 INV2 $T=1019900 1011480 1 0 $X=1019900 $Y=1006060
X3562 6076 6010 1 2 INV2 $T=1032920 981240 0 180 $X=1031060 $Y=975820
X3563 1100 6277 1 2 INV2 $T=1070120 1011480 1 0 $X=1070120 $Y=1006060
X3564 1216 6130 1 2 INV2 $T=1076940 971160 0 0 $X=1076940 $Y=970780
X3565 6488 6412 1 2 INV2 $T=1112900 1001400 1 0 $X=1112900 $Y=995980
X3566 2540 2539 1 2 BUF2 $T=407340 1001400 0 0 $X=407340 $Y=1001020
X3567 2726 2682 1 2 BUF2 $T=438340 930840 1 0 $X=438340 $Y=925420
X3568 719 4498 1 2 BUF2 $T=758260 910680 1 0 $X=758260 $Y=905260
X3569 4894 4848 1 2 BUF2 $T=819640 1021560 1 0 $X=819640 $Y=1016140
X3570 883 5065 1 2 BUF2 $T=851260 1061880 0 0 $X=851260 $Y=1061500
X3571 4703 5176 1 2 BUF2 $T=871720 961080 0 0 $X=871720 $Y=960700
X3572 5176 5598 1 2 BUF2 $T=943640 1011480 0 0 $X=943640 $Y=1011100
X3573 5990 6007 1 2 BUF2 $T=1016180 930840 0 0 $X=1016180 $Y=930460
X3574 958 1142 1 2 BUF2 $T=1019280 930840 0 0 $X=1019280 $Y=930460
X3575 6024 6064 1 2 BUF2 $T=1030440 1001400 1 0 $X=1030440 $Y=995980
X3576 970 6227 1 2 BUF2 $T=1059580 1041720 1 0 $X=1059580 $Y=1036300
X3577 1350 1 1315 1334 2 1333 ND3 $T=228160 1031640 0 180 $X=225680 $Y=1026220
X3578 1393 1 1378 1324 2 11 ND3 $T=234980 1031640 0 180 $X=232500 $Y=1026220
X3579 1446 1 1386 1360 2 1389 ND3 $T=242420 1031640 1 180 $X=239940 $Y=1031260
X3580 1397 1 1410 1491 2 1452 ND3 $T=248000 1031640 0 180 $X=245520 $Y=1026220
X3581 1572 1 1417 1500 2 1538 ND3 $T=261020 1031640 0 180 $X=258540 $Y=1026220
X3582 1596 1 37 1516 2 1576 ND3 $T=264120 940920 1 180 $X=261640 $Y=940540
X3583 1654 1 56 1642 2 1550 ND3 $T=276520 930840 0 180 $X=274040 $Y=925420
X3584 1715 1 56 1659 2 1695 ND3 $T=280860 961080 0 180 $X=278380 $Y=955660
X3585 1733 1 1609 1687 2 41 ND3 $T=283340 1021560 0 180 $X=280860 $Y=1016140
X3586 1702 1 53 1730 2 1576 ND3 $T=282100 951000 0 0 $X=282100 $Y=950620
X3587 1724 1 1630 1711 2 1389 ND3 $T=284580 1021560 0 0 $X=284580 $Y=1021180
X3588 1937 1 85 88 2 1941 ND3 $T=313720 1082040 1 180 $X=311240 $Y=1081660
X3589 1965 1 1913 1938 2 1820 ND3 $T=315580 1031640 1 180 $X=313100 $Y=1031260
X3590 1955 1 1943 1947 2 1695 ND3 $T=316820 961080 1 180 $X=314340 $Y=960700
X3591 1950 1 1717 1951 2 1689 ND3 $T=316820 1051800 0 180 $X=314340 $Y=1046380
X3592 1904 1 1717 1958 2 1754 ND3 $T=314960 1041720 1 0 $X=314960 $Y=1036300
X3593 1959 1 1695 1960 2 1902 ND3 $T=319300 951000 0 180 $X=316820 $Y=945580
X3594 1991 1 98 1996 2 122 ND3 $T=323640 910680 0 0 $X=323640 $Y=910300
X3595 1984 1 1808 1915 2 1689 ND3 $T=323640 1041720 0 0 $X=323640 $Y=1041340
X3596 2025 1 1808 2023 2 119 ND3 $T=329220 1031640 1 0 $X=329220 $Y=1026220
X3597 2009 1 133 131 2 54 ND3 $T=333560 900600 1 180 $X=331080 $Y=900220
X3598 2006 1 2055 2031 2 54 ND3 $T=334180 910680 1 180 $X=331700 $Y=910300
X3599 2041 1 136 2066 2 2055 ND3 $T=336040 920760 0 180 $X=333560 $Y=915340
X3600 2040 1 136 2091 2 133 ND3 $T=334180 910680 0 0 $X=334180 $Y=910300
X3601 2046 1 2071 2075 2 101 ND3 $T=334180 951000 1 0 $X=334180 $Y=945580
X3602 2085 1 1906 2124 2 2071 ND3 $T=339760 940920 1 0 $X=339760 $Y=935500
X3603 2065 1 2055 2117 2 2071 ND3 $T=343480 940920 0 0 $X=343480 $Y=940540
X3604 214 1 2435 215 2 2434 ND3 $T=393700 1082040 1 180 $X=391220 $Y=1081660
X3605 2500 1 2466 2495 2 2436 ND3 $T=402380 1071960 1 180 $X=399900 $Y=1071580
X3606 2529 1 2482 2512 2 2428 ND3 $T=406100 1071960 0 180 $X=403620 $Y=1066540
X3607 2563 1 2560 2553 2 2455 ND3 $T=411680 1071960 0 180 $X=409200 $Y=1066540
X3608 2569 1 2574 2596 2 2581 ND3 $T=412300 981240 0 0 $X=412300 $Y=980860
X3609 2621 1 2531 2610 2 2566 ND3 $T=420360 1001400 1 180 $X=417880 $Y=1001020
X3610 2681 1 2554 2669 2 2643 ND3 $T=429040 1001400 1 180 $X=426560 $Y=1001020
X3611 2696 1 2673 2701 2 255 ND3 $T=432140 1071960 1 0 $X=432140 $Y=1066540
X3612 2692 1 2716 2723 2 2724 ND3 $T=435860 1071960 1 0 $X=435860 $Y=1066540
X3613 2783 1 2761 2789 2 2763 ND3 $T=447020 1071960 0 180 $X=444540 $Y=1066540
X3614 2784 1 2737 2796 2 2775 ND3 $T=448880 981240 0 180 $X=446400 $Y=975820
X3615 2803 1 2801 2808 2 2770 ND3 $T=451360 951000 0 0 $X=451360 $Y=950620
X3616 2835 1 2826 2839 2 2802 ND3 $T=457560 951000 0 180 $X=455080 $Y=945580
X3617 2846 1 2714 2849 2 2854 ND3 $T=458800 1041720 1 0 $X=458800 $Y=1036300
X3618 2856 1 2779 2859 2 2855 ND3 $T=460660 1051800 1 0 $X=460660 $Y=1046380
X3619 2882 1 2815 2886 2 2891 ND3 $T=465620 991320 1 0 $X=465620 $Y=985900
X3620 2840 1 2896 2900 2 2913 ND3 $T=468720 1031640 1 0 $X=468720 $Y=1026220
X3621 2912 1 2919 2932 2 2874 ND3 $T=473060 920760 0 0 $X=473060 $Y=920380
X3622 2921 1 2924 2928 2 2866 ND3 $T=473680 920760 1 0 $X=473680 $Y=915340
X3623 2939 1 2937 2931 2 2927 ND3 $T=477400 1001400 1 180 $X=474920 $Y=1001020
X3624 2976 1 2978 2982 2 2824 ND3 $T=482360 951000 1 0 $X=482360 $Y=945580
X3625 3054 1 2995 3049 2 3019 ND3 $T=495380 981240 1 180 $X=492900 $Y=980860
X3626 3044 1 3007 3039 2 3025 ND3 $T=496000 951000 0 180 $X=493520 $Y=945580
X3627 356 1 3155 3158 2 3055 ND3 $T=516460 1051800 0 0 $X=516460 $Y=1051420
X3628 359 1 3163 3159 2 3041 ND3 $T=519560 1071960 0 180 $X=517080 $Y=1066540
X3629 367 1 3197 3221 2 2980 ND3 $T=527620 1071960 0 0 $X=527620 $Y=1071580
X3630 386 1 3270 3266 2 3035 ND3 $T=538780 1061880 1 180 $X=536300 $Y=1061500
X3631 3268 1 3208 3287 2 3097 ND3 $T=539400 1031640 0 0 $X=539400 $Y=1031260
X3632 400 1 3304 3323 2 3075 ND3 $T=546220 1041720 1 0 $X=546220 $Y=1036300
X3633 422 1 3386 3395 2 2879 ND3 $T=559240 1061880 0 180 $X=556760 $Y=1056460
X3634 3387 1 3388 3392 2 423 ND3 $T=558000 1082040 0 0 $X=558000 $Y=1081660
X3635 433 1 3429 3424 2 426 ND3 $T=566060 1082040 0 180 $X=563580 $Y=1076620
X3636 3454 1 3483 3486 2 3089 ND3 $T=574740 1021560 1 0 $X=574740 $Y=1016140
X3637 3445 1 3494 3495 2 3129 ND3 $T=577840 1021560 0 0 $X=577840 $Y=1021180
X3638 3436 1 3512 3517 2 2968 ND3 $T=582180 1061880 0 0 $X=582180 $Y=1061500
X3639 3699 1 3700 3713 2 3688 ND3 $T=619380 1051800 1 180 $X=616900 $Y=1051420
X3640 3709 1 3678 3701 2 520 ND3 $T=619380 1061880 0 180 $X=616900 $Y=1056460
X3641 3718 1 3664 3725 2 3675 ND3 $T=621240 1051800 0 180 $X=618760 $Y=1046380
X3642 3737 1 3731 3721 2 530 ND3 $T=624340 1061880 1 180 $X=621860 $Y=1061500
X3643 3840 1 3843 3859 2 566 ND3 $T=645420 1051800 1 0 $X=645420 $Y=1046380
X3644 3888 1 3897 3875 2 583 ND3 $T=655960 1051800 0 0 $X=655960 $Y=1051420
X3645 3325 1 3803 3937 2 3946 ND3 $T=662780 971160 0 0 $X=662780 $Y=970780
X3646 3948 1 3911 3964 2 3944 ND3 $T=664640 1041720 0 0 $X=664640 $Y=1041340
X3647 3509 1 3966 3970 2 3976 ND3 $T=666500 961080 0 0 $X=666500 $Y=960700
X3648 3449 1 3955 3989 2 3995 ND3 $T=668980 961080 0 0 $X=668980 $Y=960700
X3649 3463 1 3826 3990 2 3996 ND3 $T=668980 971160 1 0 $X=668980 $Y=965740
X3650 3272 1 3777 3991 2 3997 ND3 $T=668980 971160 0 0 $X=668980 $Y=970780
X3651 3471 1 4032 4020 2 4047 ND3 $T=677040 961080 1 0 $X=677040 $Y=955660
X3652 3295 1 4018 4023 2 4050 ND3 $T=678280 961080 0 0 $X=678280 $Y=960700
X3653 4057 1 4065 4081 2 4079 ND3 $T=682620 1041720 0 0 $X=682620 $Y=1041340
X3654 4098 1 4091 4089 2 637 ND3 $T=688820 1051800 0 180 $X=686340 $Y=1046380
X3655 3470 1 4175 4049 2 4190 ND3 $T=700600 951000 0 0 $X=700600 $Y=950620
X3656 4170 1 4181 4167 2 653 ND3 $T=703080 1051800 1 180 $X=700600 $Y=1051420
X3657 3224 1 4256 4011 2 4264 ND3 $T=716100 971160 0 0 $X=716100 $Y=970780
X3658 4290 1 4289 4279 2 679 ND3 $T=724160 1031640 1 180 $X=721680 $Y=1031260
X3659 3406 1 4296 4299 2 4304 ND3 $T=723540 951000 1 0 $X=723540 $Y=945580
X3660 4284 1 4311 685 2 4021 ND3 $T=725400 920760 0 0 $X=725400 $Y=920380
X3661 4275 1 4326 4339 2 692 ND3 $T=726640 1061880 1 0 $X=726640 $Y=1056460
X3662 4348 1 4355 4367 2 4329 ND3 $T=730980 1051800 0 0 $X=730980 $Y=1051420
X3663 4346 1 4363 4360 2 4349 ND3 $T=732220 1061880 0 0 $X=732220 $Y=1061500
X3664 769 1 4053 4624 2 4638 ND3 $T=780580 1001400 0 0 $X=780580 $Y=1001020
X3665 772 1 4272 4591 2 4652 ND3 $T=781820 1041720 0 0 $X=781820 $Y=1041340
X3666 773 1 4166 4647 2 4657 ND3 $T=783060 1051800 0 0 $X=783060 $Y=1051420
X3667 4664 1 4677 787 2 4608 ND3 $T=786780 910680 0 180 $X=784300 $Y=905260
X3668 780 1 4336 4634 2 4672 ND3 $T=785540 1051800 0 0 $X=785540 $Y=1051420
X3669 4679 1 4682 4675 2 4564 ND3 $T=789880 1011480 1 180 $X=787400 $Y=1011100
X3670 4697 1 4693 4685 2 4574 ND3 $T=791740 991320 1 180 $X=789260 $Y=990940
X3671 795 1 4093 4699 2 4694 ND3 $T=793600 1031640 0 180 $X=791120 $Y=1026220
X3672 790 1 4361 4680 2 4716 ND3 $T=791120 1041720 1 0 $X=791120 $Y=1036300
X3673 4711 1 4714 4702 2 4586 ND3 $T=794840 971160 0 180 $X=792360 $Y=965740
X3674 4710 1 4715 4720 2 4551 ND3 $T=792980 981240 0 0 $X=792980 $Y=980860
X3675 801 1 4362 4700 2 4735 ND3 $T=794220 1051800 0 0 $X=794220 $Y=1051420
X3676 811 1 3735 4661 2 4749 ND3 $T=794840 1051800 1 0 $X=794840 $Y=1046380
X3677 4755 1 4746 4736 2 4561 ND3 $T=798560 981240 1 180 $X=796080 $Y=980860
X3678 4698 1 4739 4738 2 4550 ND3 $T=796080 1011480 1 0 $X=796080 $Y=1006060
X3679 807 1 3690 4688 2 4752 ND3 $T=796080 1041720 0 0 $X=796080 $Y=1041340
X3680 4756 1 4747 4706 2 4558 ND3 $T=798560 1061880 0 180 $X=796080 $Y=1056460
X3681 4753 1 4748 4741 2 4559 ND3 $T=798560 1071960 1 180 $X=796080 $Y=1071580
X3682 4737 1 4740 4743 2 4573 ND3 $T=796080 1082040 1 0 $X=796080 $Y=1076620
X3683 812 1 3968 4613 2 4765 ND3 $T=798560 1011480 1 0 $X=798560 $Y=1006060
X3684 4824 1 4808 4788 2 4590 ND3 $T=807860 981240 0 180 $X=805380 $Y=975820
X3685 819 1 3881 4650 2 4826 ND3 $T=806620 1021560 0 0 $X=806620 $Y=1021180
X3686 4616 1 4817 4825 2 4821 ND3 $T=807240 940920 1 0 $X=807240 $Y=935500
X3687 4678 1 4828 4838 2 4842 ND3 $T=809100 940920 0 0 $X=809100 $Y=940540
X3688 820 1 3736 4726 2 4843 ND3 $T=809100 1021560 0 0 $X=809100 $Y=1021180
X3689 4598 1 4831 4868 2 4841 ND3 $T=810340 961080 0 0 $X=810340 $Y=960700
X3690 824 1 3715 4663 2 4858 ND3 $T=812200 1051800 0 0 $X=812200 $Y=1051420
X3691 4728 1 4887 4893 2 4827 ND3 $T=817780 951000 0 0 $X=817780 $Y=950620
X3692 4572 1 4889 4905 2 4866 ND3 $T=817780 971160 1 0 $X=817780 $Y=965740
X3693 4962 1 4983 4984 2 4987 ND3 $T=836380 981240 0 0 $X=836380 $Y=980860
X3694 4964 1 4994 4998 2 4993 ND3 $T=839480 991320 1 0 $X=839480 $Y=985900
X3695 5028 1 5039 5057 2 5062 ND3 $T=848780 991320 1 0 $X=848780 $Y=985900
X3696 5146 1 5082 5125 2 5135 ND3 $T=861800 1071960 1 0 $X=861800 $Y=1066540
X3697 5129 1 5141 5144 2 5148 ND3 $T=863660 991320 0 0 $X=863660 $Y=990940
X3698 5158 1 5126 5168 2 5181 ND3 $T=866760 1082040 1 0 $X=866760 $Y=1076620
X3699 5172 1 5116 5166 2 5159 ND3 $T=869860 991320 1 180 $X=867380 $Y=990940
X3700 5205 1 5180 5206 2 5191 ND3 $T=874820 991320 1 180 $X=872340 $Y=990940
X3701 5161 1 5059 5198 2 5210 ND3 $T=872960 1061880 0 0 $X=872960 $Y=1061500
X3702 5239 1 5227 5231 2 5220 ND3 $T=880400 991320 0 180 $X=877920 $Y=985900
X3703 5342 1 5343 5357 2 5324 ND3 $T=897140 971160 0 0 $X=897140 $Y=970780
X3704 5350 1 5360 5369 2 5363 ND3 $T=897760 961080 1 0 $X=897760 $Y=955660
X3705 5356 1 5400 5402 2 5294 ND3 $T=906440 961080 1 0 $X=906440 $Y=955660
X3706 5378 1 5401 5403 2 5215 ND3 $T=906440 991320 0 0 $X=906440 $Y=990940
X3707 5322 1 5416 5422 2 5379 ND3 $T=912640 971160 0 0 $X=912640 $Y=970780
X3708 5456 1 981 4732 2 5471 ND3 $T=920700 1051800 1 0 $X=920700 $Y=1046380
X3709 5459 1 5466 4723 2 5477 ND3 $T=921320 1061880 0 0 $X=921320 $Y=1061500
X3710 5482 1 989 4758 2 5495 ND3 $T=923800 1071960 1 0 $X=923800 $Y=1066540
X3711 5530 1 1005 4690 2 1001 ND3 $T=933100 1082040 1 180 $X=930620 $Y=1081660
X3712 5531 1 5525 4885 2 5519 ND3 $T=933720 951000 0 180 $X=931240 $Y=945580
X3713 5541 1 5546 4878 2 5552 ND3 $T=934960 940920 1 0 $X=934960 $Y=935500
X3714 5574 1 1020 4790 2 5586 ND3 $T=939920 1041720 0 0 $X=939920 $Y=1041340
X3715 5585 1 5591 5026 2 5601 ND3 $T=941780 951000 0 0 $X=941780 $Y=950620
X3716 5588 1 5606 4907 2 5614 ND3 $T=944880 981240 0 0 $X=944880 $Y=980860
X3717 5567 1 5611 4869 2 5620 ND3 $T=945500 1011480 1 0 $X=945500 $Y=1006060
X3718 5566 1 5621 4705 2 5632 ND3 $T=946740 1011480 0 0 $X=946740 $Y=1011100
X3719 5642 1 5637 5475 2 5625 ND3 $T=950460 961080 0 180 $X=947980 $Y=955660
X3720 5651 1 5661 5169 2 1034 ND3 $T=952320 1071960 1 0 $X=952320 $Y=1066540
X3721 5668 1 1038 5174 2 5690 ND3 $T=956040 1031640 1 0 $X=956040 $Y=1026220
X3722 5698 1 5670 5212 2 5708 ND3 $T=959760 1011480 1 0 $X=959760 $Y=1006060
X3723 5649 1 1044 5131 2 5713 ND3 $T=960380 1061880 0 0 $X=960380 $Y=1061500
X3724 5701 1 5695 5052 2 5714 ND3 $T=960380 1071960 1 0 $X=960380 $Y=1066540
X3725 5712 1 1049 5058 2 5720 ND3 $T=962240 1021560 0 0 $X=962240 $Y=1021180
X3726 5744 1 5742 5374 2 5735 ND3 $T=969060 971160 0 180 $X=966580 $Y=965740
X3727 5709 1 1060 5228 2 5745 ND3 $T=966580 1051800 1 0 $X=966580 $Y=1046380
X3728 5758 1 5706 5461 2 5752 ND3 $T=968440 991320 0 0 $X=968440 $Y=990940
X3729 5751 1 5693 5494 2 5762 ND3 $T=970300 971160 0 0 $X=970300 $Y=970780
X3730 5780 1 5771 5474 2 5787 ND3 $T=975880 940920 0 0 $X=975880 $Y=940540
X3731 1324 1323 1334 2 1 ND2S $T=224440 1021560 1 180 $X=222580 $Y=1021180
X3732 1333 1319 1350 2 1 ND2S $T=225680 1021560 0 0 $X=225680 $Y=1021180
X3733 1338 1346 1333 2 1 ND2S $T=230020 1021560 1 180 $X=228160 $Y=1021180
X3734 11 1341 1378 2 1 ND2S $T=230020 1021560 0 0 $X=230020 $Y=1021180
X3735 1389 1383 1350 2 1 ND2S $T=233740 1021560 1 180 $X=231880 $Y=1021180
X3736 18 1434 1403 2 1 ND2S $T=238700 1031640 1 180 $X=236840 $Y=1031260
X3737 1452 1401 1386 2 1 ND2S $T=238700 1021560 0 0 $X=238700 $Y=1021180
X3738 1452 1408 1397 2 1 ND2S $T=242420 1031640 1 0 $X=242420 $Y=1026220
X3739 1389 1453 1386 2 1 ND2S $T=244280 1031640 1 180 $X=242420 $Y=1031260
X3740 1500 1478 1491 2 1 ND2S $T=249860 1031640 0 180 $X=248000 $Y=1026220
X3741 31 1474 25 2 1 ND2S $T=251100 910680 0 180 $X=249240 $Y=905260
X3742 1333 1504 1397 2 1 ND2S $T=251100 1031640 1 180 $X=249240 $Y=1031260
X3743 27 1507 25 2 1 ND2S $T=251100 910680 1 0 $X=251100 $Y=905260
X3744 29 1512 1397 2 1 ND2S $T=252960 1011480 0 180 $X=251100 $Y=1006060
X3745 1538 1495 1417 2 1 ND2S $T=251100 1021560 0 0 $X=251100 $Y=1021180
X3746 25 30 32 2 1 ND2S $T=252960 900600 0 0 $X=252960 $Y=900220
X3747 1389 1510 1397 2 1 ND2S $T=254820 1031640 1 180 $X=252960 $Y=1031260
X3748 27 1523 37 2 1 ND2S $T=256060 940920 0 0 $X=256060 $Y=940540
X3749 34 1522 1554 2 1 ND2S $T=256060 1011480 0 0 $X=256060 $Y=1011100
X3750 31 1545 37 2 1 ND2S $T=256680 940920 1 0 $X=256680 $Y=935500
X3751 14 1553 1541 2 1 ND2S $T=258540 1021560 0 180 $X=256680 $Y=1016140
X3752 34 1534 1378 2 1 ND2S $T=258540 1031640 1 180 $X=256680 $Y=1031260
X3753 37 1540 32 2 1 ND2S $T=258540 920760 1 0 $X=258540 $Y=915340
X3754 1570 1558 1545 2 1 ND2S $T=260400 940920 1 180 $X=258540 $Y=940540
X3755 1576 1570 43 2 1 ND2S $T=261640 951000 0 0 $X=261640 $Y=950620
X3756 41 1438 1608 2 1 ND2S $T=263500 1011480 0 0 $X=263500 $Y=1011100
X3757 1550 1617 43 2 1 ND2S $T=267220 920760 1 180 $X=265360 $Y=920380
X3758 46 1511 1544 2 1 ND2S $T=265360 1031640 1 0 $X=265360 $Y=1026220
X3759 40 1567 1403 2 1 ND2S $T=265980 1041720 1 0 $X=265980 $Y=1036300
X3760 1452 1620 1544 2 1 ND2S $T=269080 1031640 1 180 $X=267220 $Y=1031260
X3761 1538 1592 1586 2 1 ND2S $T=267220 1041720 0 0 $X=267220 $Y=1041340
X3762 53 1650 32 2 1 ND2S $T=270940 951000 0 180 $X=269080 $Y=945580
X3763 1677 1548 1644 2 1 ND2S $T=272180 1041720 1 180 $X=270320 $Y=1041340
X3764 41 1652 1378 2 1 ND2S $T=272800 1031640 1 180 $X=270940 $Y=1031260
X3765 1567 1664 1652 2 1 ND2S $T=270940 1041720 1 0 $X=270940 $Y=1036300
X3766 54 1619 53 2 1 ND2S $T=272180 920760 0 0 $X=272180 $Y=920380
X3767 1672 1647 1642 2 1 ND2S $T=274040 940920 0 180 $X=272180 $Y=935500
X3768 1615 1601 53 2 1 ND2S $T=272180 951000 0 0 $X=272180 $Y=950620
X3769 1678 1656 1662 2 1 ND2S $T=272180 961080 1 0 $X=272180 $Y=955660
X3770 40 1566 1644 2 1 ND2S $T=272180 1011480 0 0 $X=272180 $Y=1011100
X3771 1538 1661 1644 2 1 ND2S $T=274040 1041720 1 180 $X=272180 $Y=1041340
X3772 1550 1632 60 2 1 ND2S $T=274040 920760 0 0 $X=274040 $Y=920380
X3773 1681 1672 1632 2 1 ND2S $T=275900 940920 0 180 $X=274040 $Y=935500
X3774 1333 1684 1417 2 1 ND2S $T=275900 1031640 1 180 $X=274040 $Y=1031260
X3775 1677 1671 1586 2 1 ND2S $T=275900 1041720 1 180 $X=274040 $Y=1041340
X3776 1659 1666 1678 2 1 ND2S $T=274660 951000 0 0 $X=274660 $Y=950620
X3777 1689 1676 1417 2 1 ND2S $T=277760 1051800 0 180 $X=275900 $Y=1046380
X3778 1695 1681 56 2 1 ND2S $T=278380 940920 0 180 $X=276520 $Y=935500
X3779 1576 1697 60 2 1 ND2S $T=279620 940920 1 180 $X=277760 $Y=940540
X3780 1687 1692 1690 2 1 ND2S $T=279620 1021560 0 180 $X=277760 $Y=1016140
X3781 1688 1686 1664 2 1 ND2S $T=279000 1041720 1 0 $X=279000 $Y=1036300
X3782 41 1707 1403 2 1 ND2S $T=283340 1031640 1 0 $X=283340 $Y=1026220
X3783 1389 1764 1630 2 1 ND2S $T=288300 1021560 0 180 $X=286440 $Y=1016140
X3784 1749 1758 1717 2 1 ND2S $T=287680 1041720 0 0 $X=287680 $Y=1041340
X3785 1754 1769 1630 2 1 ND2S $T=290160 1041720 0 180 $X=288300 $Y=1036300
X3786 46 1776 1800 2 1 ND2S $T=292640 1031640 0 0 $X=292640 $Y=1031260
X3787 32 1806 67 2 1 ND2S $T=295120 951000 0 0 $X=295120 $Y=950620
X3788 1615 1829 67 2 1 ND2S $T=297600 961080 0 180 $X=295740 $Y=955660
X3789 46 1768 1674 2 1 ND2S $T=296980 1031640 0 0 $X=296980 $Y=1031260
X3790 1803 1835 1819 2 1 ND2S $T=299460 961080 0 180 $X=297600 $Y=955660
X3791 1835 1824 1856 2 1 ND2S $T=298840 961080 0 0 $X=298840 $Y=960700
X3792 1754 1847 1586 2 1 ND2S $T=301320 1041720 0 180 $X=299460 $Y=1036300
X3793 1689 1850 1586 2 1 ND2S $T=301320 1041720 1 180 $X=299460 $Y=1041340
X3794 79 1821 1808 2 1 ND2S $T=303800 1051800 1 0 $X=303800 $Y=1046380
X3795 1894 1892 1714 2 1 ND2S $T=307520 930840 1 180 $X=305660 $Y=930460
X3796 1894 1889 89 2 1 ND2S $T=306280 920760 0 0 $X=306280 $Y=920380
X3797 1892 1873 1866 2 1 ND2S $T=306280 940920 0 0 $X=306280 $Y=940540
X3798 1820 1898 1800 2 1 ND2S $T=308140 1031640 1 180 $X=306280 $Y=1031260
X3799 1889 1859 1905 2 1 ND2S $T=306900 920760 1 0 $X=306900 $Y=915340
X3800 1902 1828 90 2 1 ND2S $T=307520 951000 1 0 $X=307520 $Y=945580
X3801 90 1762 1906 2 1 ND2S $T=310000 930840 1 180 $X=308140 $Y=930460
X3802 1906 1823 95 2 1 ND2S $T=308140 940920 1 0 $X=308140 $Y=935500
X3803 1902 1777 95 2 1 ND2S $T=308140 951000 0 0 $X=308140 $Y=950620
X3804 1820 1827 1913 2 1 ND2S $T=308140 1031640 0 0 $X=308140 $Y=1031260
X3805 94 1771 98 2 1 ND2S $T=310000 930840 0 0 $X=310000 $Y=930460
X3806 1902 1900 94 2 1 ND2S $T=310000 951000 1 0 $X=310000 $Y=945580
X3807 1749 1914 1913 2 1 ND2S $T=310000 1031640 0 0 $X=310000 $Y=1031260
X3808 1928 1862 95 2 1 ND2S $T=313100 961080 0 180 $X=311240 $Y=955660
X3809 1928 1858 104 2 1 ND2S $T=313100 930840 1 0 $X=313100 $Y=925420
X3810 1938 1954 1958 2 1 ND2S $T=315580 1031640 0 0 $X=315580 $Y=1031260
X3811 1947 1969 1963 2 1 ND2S $T=316820 971160 0 0 $X=316820 $Y=970780
X3812 1754 1970 1717 2 1 ND2S $T=319300 1041720 0 180 $X=317440 $Y=1036300
X3813 1749 1926 1800 2 1 ND2S $T=318680 1031640 1 0 $X=318680 $Y=1026220
X3814 1963 1961 1973 2 1 ND2S $T=319300 971160 1 0 $X=319300 $Y=965740
X3815 1965 1983 1879 2 1 ND2S $T=320540 1031640 0 0 $X=320540 $Y=1031260
X3816 117 1937 1953 2 1 ND2S $T=320540 1082040 1 0 $X=320540 $Y=1076620
X3817 1689 1962 1717 2 1 ND2S $T=321160 1051800 1 0 $X=321160 $Y=1046380
X3818 1615 1982 1928 2 1 ND2S $T=321780 961080 1 0 $X=321780 $Y=955660
X3819 1992 1993 1994 2 1 ND2S $T=324260 961080 0 0 $X=324260 $Y=960700
X3820 129 2016 1800 2 1 ND2S $T=329220 1021560 1 180 $X=327360 $Y=1021180
X3821 129 1995 1808 2 1 ND2S $T=329220 1041720 0 180 $X=327360 $Y=1036300
X3822 119 2029 1808 2 1 ND2S $T=331080 1031640 1 180 $X=329220 $Y=1031260
X3823 1983 2049 2023 2 1 ND2S $T=332940 1031640 1 180 $X=331080 $Y=1031260
X3824 1996 2051 2066 2 1 ND2S $T=331700 920760 1 0 $X=331700 $Y=915340
X3825 1928 2059 136 2 1 ND2S $T=332940 920760 0 0 $X=332940 $Y=920380
X3826 133 2082 136 2 1 ND2S $T=336040 900600 1 180 $X=334180 $Y=900220
X3827 139 2076 133 2 1 ND2S $T=336660 930840 0 180 $X=334800 $Y=925420
X3828 2031 2099 2091 2 1 ND2S $T=337900 920760 0 180 $X=336040 $Y=915340
X3829 140 2104 2081 2 1 ND2S $T=337900 1061880 1 180 $X=336040 $Y=1061500
X3830 135 2100 133 2 1 ND2S $T=338520 920760 1 180 $X=336660 $Y=920380
X3831 2055 2095 136 2 1 ND2S $T=339760 910680 1 180 $X=337900 $Y=910300
X3832 135 2112 2055 2 1 ND2S $T=337900 930840 1 0 $X=337900 $Y=925420
X3833 141 2110 2081 2 1 ND2S $T=339760 1071960 1 180 $X=337900 $Y=1071580
X3834 2117 2116 2086 2 1 ND2S $T=341620 951000 0 180 $X=339760 $Y=945580
X3835 148 1957 2137 2 1 ND2S $T=339760 1082040 0 0 $X=339760 $Y=1081660
X3836 129 2121 1913 2 1 ND2S $T=343480 1031640 0 180 $X=341620 $Y=1026220
X3837 2071 2150 2055 2 1 ND2S $T=345340 940920 0 180 $X=343480 $Y=935500
X3838 119 2159 1912 2 1 ND2S $T=347200 1021560 1 180 $X=345340 $Y=1021180
X3839 138 2135 158 2 1 ND2S $T=345340 1082040 1 0 $X=345340 $Y=1076620
X3840 164 2177 1807 2 1 ND2S $T=352160 1001400 1 180 $X=350300 $Y=1001020
X3841 95 2136 166 2 1 ND2S $T=350920 940920 0 0 $X=350920 $Y=940540
X3842 2197 2198 2191 2 1 ND2S $T=354020 1031640 0 180 $X=352160 $Y=1026220
X3843 94 2213 177 2 1 ND2S $T=360220 951000 1 0 $X=360220 $Y=945580
X3844 95 2209 177 2 1 ND2S $T=360840 940920 1 0 $X=360840 $Y=935500
X3845 2269 2311 2238 2 1 ND2S $T=372000 951000 0 180 $X=370140 $Y=945580
X3846 2311 2271 2265 2 1 ND2S $T=372000 951000 1 180 $X=370140 $Y=950620
X3847 2262 2319 2269 2 1 ND2S $T=373240 940920 1 180 $X=371380 $Y=940540
X3848 104 2316 166 2 1 ND2S $T=372000 920760 0 0 $X=372000 $Y=920380
X3849 2361 2318 2351 2 1 ND2S $T=375720 930840 0 0 $X=375720 $Y=930460
X3850 2228 2361 2363 2 1 ND2S $T=377580 930840 0 0 $X=377580 $Y=930460
X3851 2228 2378 199 2 1 ND2S $T=382540 920760 0 0 $X=382540 $Y=920380
X3852 2378 2371 2400 2 1 ND2S $T=384400 930840 0 0 $X=384400 $Y=930460
X3853 2431 2425 2319 2 1 ND2S $T=390600 930840 0 0 $X=390600 $Y=930460
X3854 2319 2448 213 2 1 ND2S $T=393700 940920 0 180 $X=391840 $Y=935500
X3855 2463 2431 213 2 1 ND2S $T=394320 930840 1 180 $X=392460 $Y=930460
X3856 217 2503 2463 2 1 ND2S $T=400520 940920 0 180 $X=398660 $Y=935500
X3857 2503 2489 221 2 1 ND2S $T=402380 940920 0 180 $X=400520 $Y=935500
X3858 2535 2529 2528 2 1 ND2S $T=406100 1071960 1 0 $X=406100 $Y=1066540
X3859 2535 2500 2502 2 1 ND2S $T=406720 1071960 0 0 $X=406720 $Y=1071580
X3860 2535 2563 2571 2 1 ND2S $T=415400 1071960 0 0 $X=415400 $Y=1071580
X3861 2634 2569 2639 2 1 ND2S $T=420980 1001400 1 0 $X=420980 $Y=995980
X3862 2634 2621 2611 2 1 ND2S $T=421600 1001400 0 0 $X=421600 $Y=1001020
X3863 2634 2681 2652 2 1 ND2S $T=427180 1011480 1 0 $X=427180 $Y=1006060
X3864 2535 2692 2647 2 1 ND2S $T=430280 1071960 1 180 $X=428420 $Y=1071580
X3865 2535 2696 2620 2 1 ND2S $T=430900 1071960 0 180 $X=429040 $Y=1066540
X3866 2759 2691 2778 2 1 ND2S $T=444540 1001400 0 0 $X=444540 $Y=1001020
X3867 2793 2783 2772 2 1 ND2S $T=447020 1061880 0 180 $X=445160 $Y=1056460
X3868 2786 2784 2776 2 1 ND2S $T=448260 981240 1 180 $X=446400 $Y=980860
X3869 2786 2803 2811 2 1 ND2S $T=451980 961080 1 0 $X=451980 $Y=955660
X3870 2786 2835 2797 2 1 ND2S $T=456940 951000 0 0 $X=456940 $Y=950620
X3871 2793 2846 2834 2 1 ND2S $T=458800 1041720 0 180 $X=456940 $Y=1036300
X3872 2793 2840 2809 2 1 ND2S $T=459420 1021560 1 180 $X=457560 $Y=1021180
X3873 2793 2856 2843 2 1 ND2S $T=460660 1051800 0 180 $X=458800 $Y=1046380
X3874 2786 2882 2864 2 1 ND2S $T=465620 991320 0 180 $X=463760 $Y=985900
X3875 302 2912 2862 2 1 ND2S $T=471820 920760 0 180 $X=469960 $Y=915340
X3876 302 2921 2853 2 1 ND2S $T=473680 920760 0 180 $X=471820 $Y=915340
X3877 302 304 2901 2 1 ND2S $T=476160 910680 0 180 $X=474300 $Y=905260
X3878 2786 2939 2949 2 1 ND2S $T=476780 991320 1 0 $X=476780 $Y=985900
X3879 2940 2936 2954 2 1 ND2S $T=477400 940920 1 0 $X=477400 $Y=935500
X3880 314 2976 2962 2 1 ND2S $T=484220 961080 0 180 $X=482360 $Y=955660
X3881 314 3054 3018 2 1 ND2S $T=500340 981240 1 0 $X=500340 $Y=975820
X3882 314 3044 3073 2 1 ND2S $T=503440 961080 1 0 $X=503440 $Y=955660
X3883 779 4664 4648 2 1 ND2S $T=786160 910680 1 180 $X=784300 $Y=910300
X3884 4686 4679 4612 2 1 ND2S $T=789880 1001400 1 180 $X=788020 $Y=1001020
X3885 4686 4710 4617 2 1 ND2S $T=792980 981240 1 180 $X=791120 $Y=980860
X3886 4686 4698 4656 2 1 ND2S $T=792980 1011480 0 180 $X=791120 $Y=1006060
X3887 796 4737 793 2 1 ND2S $T=793600 1082040 0 180 $X=791740 $Y=1076620
X3888 4686 4697 4581 2 1 ND2S $T=792360 991320 0 0 $X=792360 $Y=990940
X3889 4686 4711 4625 2 1 ND2S $T=794840 971160 1 180 $X=792980 $Y=970780
X3890 4718 4682 4689 2 1 ND2S $T=794220 1011480 1 0 $X=794220 $Y=1006060
X3891 4718 4693 4733 2 1 ND2S $T=794840 991320 0 0 $X=794840 $Y=990940
X3892 4718 4714 4549 2 1 ND2S $T=796080 971160 0 0 $X=796080 $Y=970780
X3893 4718 4715 4514 2 1 ND2S $T=796700 991320 1 0 $X=796700 $Y=985900
X3894 4727 4756 4724 2 1 ND2S $T=798560 1061880 1 180 $X=796700 $Y=1061500
X3895 4727 4753 4605 2 1 ND2S $T=798560 1071960 0 180 $X=796700 $Y=1066540
X3896 4686 4755 4713 2 1 ND2S $T=798560 991320 1 0 $X=798560 $Y=985900
X3897 4718 4739 4784 2 1 ND2S $T=801660 1001400 0 0 $X=801660 $Y=1001020
X3898 4782 4824 4818 2 1 ND2S $T=807860 971160 0 0 $X=807860 $Y=970780
X3899 4718 4746 4839 2 1 ND2S $T=809100 981240 0 0 $X=809100 $Y=980860
X3900 4813 4808 4845 2 1 ND2S $T=810340 971160 0 0 $X=810340 $Y=970780
X3901 4871 4880 4772 2 1 ND2S $T=816540 920760 0 180 $X=814680 $Y=915340
X3902 789 4877 4874 2 1 ND2S $T=817780 920760 1 0 $X=817780 $Y=915340
X3903 4782 4962 4946 2 1 ND2S $T=833900 981240 1 180 $X=832040 $Y=980860
X3904 4924 4983 4941 2 1 ND2S $T=835760 981240 1 180 $X=833900 $Y=980860
X3905 4782 4964 4947 2 1 ND2S $T=835760 991320 0 180 $X=833900 $Y=985900
X3906 4924 4994 4972 2 1 ND2S $T=838860 991320 0 180 $X=837000 $Y=985900
X3907 5021 5028 4976 2 1 ND2S $T=844440 991320 1 180 $X=842580 $Y=990940
X3908 4924 5039 5015 2 1 ND2S $T=846300 981240 0 0 $X=846300 $Y=980860
X3909 5050 5116 5051 2 1 ND2S $T=859320 1001400 0 180 $X=857460 $Y=995980
X3910 5021 5129 5128 2 1 ND2S $T=864280 991320 0 180 $X=862420 $Y=985900
X3911 901 5158 5136 2 1 ND2S $T=865520 1082040 0 180 $X=863660 $Y=1076620
X3912 4727 5146 5154 2 1 ND2S $T=864280 1071960 1 0 $X=864280 $Y=1066540
X3913 5050 5141 5100 2 1 ND2S $T=868000 1001400 0 180 $X=866140 $Y=995980
X3914 901 5161 5123 2 1 ND2S $T=868620 1061880 1 180 $X=866760 $Y=1061500
X3915 5021 5172 5185 2 1 ND2S $T=869240 1001400 1 0 $X=869240 $Y=995980
X3916 5050 5180 5171 2 1 ND2S $T=870480 991320 0 0 $X=870480 $Y=990940
X3917 5021 5205 5202 2 1 ND2S $T=875440 991320 0 0 $X=875440 $Y=990940
X3918 916 5251 5209 2 1 ND2S $T=879780 920760 0 180 $X=877920 $Y=915340
X3919 5050 5227 5203 2 1 ND2S $T=879780 991320 1 180 $X=877920 $Y=990940
X3920 916 5240 5236 2 1 ND2S $T=881640 910680 1 180 $X=879780 $Y=910300
X3921 916 5254 5222 2 1 ND2S $T=881640 920760 0 180 $X=879780 $Y=915340
X3922 5021 5239 5259 2 1 ND2S $T=881640 991320 1 0 $X=881640 $Y=985900
X3923 835 5257 5299 2 1 ND2S $T=884120 920760 0 0 $X=884120 $Y=920380
X3924 835 5278 933 2 1 ND2S $T=887220 900600 0 0 $X=887220 $Y=900220
X3925 835 5279 5302 2 1 ND2S $T=887220 910680 1 0 $X=887220 $Y=905260
X3926 835 5292 5311 2 1 ND2S $T=888460 920760 1 0 $X=888460 $Y=915340
X3927 947 5271 5370 2 1 ND2S $T=899620 920760 1 0 $X=899620 $Y=915340
X3928 947 5303 5380 2 1 ND2S $T=900860 910680 0 0 $X=900860 $Y=910300
X3929 947 5267 5305 2 1 ND2S $T=901480 910680 1 0 $X=901480 $Y=905260
X3930 947 5266 960 2 1 ND2S $T=903340 900600 0 0 $X=903340 $Y=900220
X3931 5429 5430 5410 2 1 ND2S $T=915120 940920 1 180 $X=913260 $Y=940540
X3932 1309 1310 1 1309 1310 1304 2 MOAI1S $T=223820 1041720 0 180 $X=220100 $Y=1036300
X3933 1304 1306 1 1304 1306 1321 2 MOAI1S $T=220100 1061880 1 0 $X=220100 $Y=1056460
X3934 1315 1319 1 1315 1319 1331 2 MOAI1S $T=221340 1031640 1 0 $X=221340 $Y=1026220
X3935 1326 1339 1 1326 1314 1317 2 MOAI1S $T=227540 991320 0 180 $X=223820 $Y=985900
X3936 1326 1345 1 1326 1330 1308 2 MOAI1S $T=228160 1001400 0 180 $X=224440 $Y=995980
X3937 1335 1332 1 1335 1332 1310 2 MOAI1S $T=228160 1041720 0 180 $X=224440 $Y=1036300
X3938 1336 1342 1 1336 1342 1361 2 MOAI1S $T=225680 1061880 1 0 $X=225680 $Y=1056460
X3939 1341 1346 1 1341 1346 1367 2 MOAI1S $T=226300 1021560 1 0 $X=226300 $Y=1016140
X3940 1326 1374 1 1326 10 1316 2 MOAI1S $T=231880 991320 0 180 $X=228160 $Y=985900
X3941 1365 1360 1 1365 1360 1332 2 MOAI1S $T=232500 1041720 0 180 $X=228780 $Y=1036300
X3942 1375 1361 1 1375 1361 1306 2 MOAI1S $T=233740 1061880 0 180 $X=230020 $Y=1056460
X3943 1369 1367 1 1369 1367 1391 2 MOAI1S $T=230640 1021560 1 0 $X=230640 $Y=1016140
X3944 1387 1391 1 1387 1391 1416 2 MOAI1S $T=233120 1011480 1 0 $X=233120 $Y=1006060
X3945 1401 1383 1 1401 1383 1369 2 MOAI1S $T=237460 1021560 1 180 $X=233740 $Y=1021180
X3946 1410 1408 1 1410 1408 1392 2 MOAI1S $T=238700 1031640 0 180 $X=234980 $Y=1026220
X3947 1429 1416 1 1429 1416 1322 2 MOAI1S $T=241180 1011480 0 180 $X=237460 $Y=1006060
X3948 1434 1438 1 1434 1438 1387 2 MOAI1S $T=242420 1011480 1 180 $X=238700 $Y=1011100
X3949 1447 1461 1 1447 1461 1309 2 MOAI1S $T=246760 1011480 1 180 $X=243040 $Y=1011100
X3950 1388 1463 1 1388 22 1477 2 MOAI1S $T=243660 1001400 1 0 $X=243660 $Y=995980
X3951 1467 1464 1 1467 1464 1342 2 MOAI1S $T=247380 1051800 0 180 $X=243660 $Y=1046380
X3952 1446 1453 1 1446 1453 1488 2 MOAI1S $T=244900 1031640 0 0 $X=244900 $Y=1031260
X3953 1380 1478 1 1380 1478 1499 2 MOAI1S $T=246140 1011480 1 0 $X=246140 $Y=1006060
X3954 1494 1489 1 1494 1489 1487 2 MOAI1S $T=251100 940920 1 180 $X=247380 $Y=940540
X3955 1495 1490 1 1495 1490 1461 2 MOAI1S $T=251100 1011480 1 180 $X=247380 $Y=1011100
X3956 1496 1501 1 1496 1501 1535 2 MOAI1S $T=248620 1051800 1 0 $X=248620 $Y=1046380
X3957 1515 1511 1 1515 1511 1439 2 MOAI1S $T=254200 1082040 0 180 $X=250480 $Y=1076620
X3958 1388 1472 1 1509 1528 1537 2 MOAI1S $T=251100 1001400 1 0 $X=251100 $Y=995980
X3959 1512 1522 1 1512 1522 1490 2 MOAI1S $T=255440 1011480 1 180 $X=251720 $Y=1011100
X3960 1514 1510 1 1514 1510 1547 2 MOAI1S $T=253580 1041720 1 0 $X=253580 $Y=1036300
X3961 1542 1540 1 1542 1540 1519 2 MOAI1S $T=258540 920760 0 180 $X=254820 $Y=915340
X3962 1400 1546 1 1400 1560 1533 2 MOAI1S $T=256060 1001400 1 0 $X=256060 $Y=995980
X3963 1553 1566 1 1553 1566 1429 2 MOAI1S $T=262260 1011480 1 180 $X=258540 $Y=1011100
X3964 1400 1577 1 1400 1591 1582 2 MOAI1S $T=260400 1001400 1 0 $X=260400 $Y=995980
X3965 44 1604 1 1574 1540 1573 2 MOAI1S $T=265360 920760 0 180 $X=261640 $Y=915340
X3966 1589 1595 1 1589 1595 1614 2 MOAI1S $T=262880 930840 1 0 $X=262880 $Y=925420
X3967 1605 1592 1 1605 1592 1563 2 MOAI1S $T=267220 1051800 1 180 $X=263500 $Y=1051420
X3968 1585 1504 1 1585 1504 1616 2 MOAI1S $T=263500 1061880 1 0 $X=263500 $Y=1056460
X3969 1639 1629 1 1639 1638 1626 2 MOAI1S $T=272180 1011480 1 180 $X=268460 $Y=1011100
X3970 1648 1627 1 1648 1627 1635 2 MOAI1S $T=273420 1051800 1 180 $X=269700 $Y=1051420
X3971 1671 1661 1 1592 1548 1627 2 MOAI1S $T=275900 1051800 0 180 $X=272180 $Y=1046380
X3972 1662 1666 1 1662 1666 1673 2 MOAI1S $T=272800 961080 0 0 $X=272800 $Y=960700
X3973 1647 1650 1 1647 1650 1663 2 MOAI1S $T=274040 940920 0 0 $X=274040 $Y=940540
X3974 46 1609 1 51 1657 1690 2 MOAI1S $T=274040 1021560 1 0 $X=274040 $Y=1016140
X3975 1669 1676 1 1669 1676 1705 2 MOAI1S $T=276520 1051800 0 0 $X=276520 $Y=1051420
X3976 1686 1684 1 1686 1684 1719 2 MOAI1S $T=278380 1051800 1 0 $X=278380 $Y=1046380
X3977 1692 1711 1 1692 1711 1712 2 MOAI1S $T=279620 1021560 0 0 $X=279620 $Y=1021180
X3978 1658 1665 1 1658 1665 1736 2 MOAI1S $T=279620 1082040 0 0 $X=279620 $Y=1081660
X3979 1744 1742 1 1744 1742 1739 2 MOAI1S $T=288300 940920 1 180 $X=284580 $Y=940540
X3980 1735 1730 1 1735 1730 1759 2 MOAI1S $T=284580 961080 1 0 $X=284580 $Y=955660
X3981 1736 1653 1 1736 1653 1780 2 MOAI1S $T=284580 1082040 0 0 $X=284580 $Y=1081660
X3982 1733 1720 1 1733 1720 1751 2 MOAI1S $T=285200 1051800 0 0 $X=285200 $Y=1051420
X3983 1724 1764 1 1724 1764 1761 2 MOAI1S $T=292020 1021560 1 180 $X=288300 $Y=1021180
X3984 1509 1767 1 1509 1782 1787 2 MOAI1S $T=288920 1001400 0 0 $X=288920 $Y=1001020
X3985 1707 1768 1 1776 1652 1785 2 MOAI1S $T=288920 1031640 0 0 $X=288920 $Y=1031260
X3986 1789 1771 1 1789 1771 1670 2 MOAI1S $T=295120 930840 1 180 $X=291400 $Y=930460
X3987 1695 67 1 1778 1746 1678 2 MOAI1S $T=295120 961080 0 180 $X=291400 $Y=955660
X3988 1828 1823 1 1762 1777 1742 2 MOAI1S $T=297600 940920 0 180 $X=293880 $Y=935500
X3989 1812 1806 1 1812 1806 1802 2 MOAI1S $T=297600 971160 0 180 $X=293880 $Y=965740
X3990 1769 1816 1 1769 1816 1841 2 MOAI1S $T=295120 1041720 1 0 $X=295120 $Y=1036300
X3991 1814 1758 1 1814 1758 1851 2 MOAI1S $T=295120 1051800 0 0 $X=295120 $Y=1051420
X3992 1811 1824 1 1811 1824 1794 2 MOAI1S $T=299460 971160 1 180 $X=295740 $Y=970780
X3993 1639 1834 1 1639 1826 1810 2 MOAI1S $T=299460 1011480 0 180 $X=295740 $Y=1006060
X3994 1876 1861 1 1845 1806 1728 2 MOAI1S $T=303180 971160 0 180 $X=299460 $Y=965740
X3995 1859 1858 1 1859 1858 1852 2 MOAI1S $T=303800 930840 0 180 $X=300080 $Y=925420
X3996 1855 1847 1 1855 1847 1885 2 MOAI1S $T=300080 1051800 1 0 $X=300080 $Y=1046380
X3997 1639 1878 1 1639 1863 1836 2 MOAI1S $T=305040 1011480 0 180 $X=301320 $Y=1006060
X3998 1862 1829 1 1862 1829 1881 2 MOAI1S $T=301940 991320 0 0 $X=301940 $Y=990940
X3999 1799 1865 1 1799 1881 1888 2 MOAI1S $T=301940 1001400 1 0 $X=301940 $Y=995980
X4000 1849 1850 1 1849 1850 1891 2 MOAI1S $T=302560 1061880 0 0 $X=302560 $Y=1061500
X4001 1872 1873 1 1872 1873 1753 2 MOAI1S $T=306900 951000 0 180 $X=303180 $Y=945580
X4002 1897 1780 1 1897 1895 1927 2 MOAI1S $T=306900 991320 1 0 $X=306900 $Y=985900
X4003 1897 1908 1 1897 1877 1924 2 MOAI1S $T=307520 991320 0 0 $X=307520 $Y=990940
X4004 1897 1499 1 1897 1922 1932 2 MOAI1S $T=308760 1001400 1 0 $X=308760 $Y=995980
X4005 101 100 1 96 81 1856 2 MOAI1S $T=313720 920760 0 180 $X=310000 $Y=915340
X4006 1943 105 1 1917 1871 1866 2 MOAI1S $T=315580 940920 1 180 $X=311860 $Y=940540
X4007 1931 1907 1 1931 1907 1797 2 MOAI1S $T=315580 971160 0 180 $X=311860 $Y=965740
X4008 1695 1928 1 1778 1880 1963 2 MOAI1S $T=313720 961080 1 0 $X=313720 $Y=955660
X4009 1950 1962 1 1950 1962 1956 2 MOAI1S $T=320540 1051800 0 180 $X=316820 $Y=1046380
X4010 112 116 1 1968 1871 1905 2 MOAI1S $T=321780 920760 0 180 $X=318060 $Y=915340
X4011 1904 1970 1 1904 1970 2036 2 MOAI1S $T=319300 1041720 0 0 $X=319300 $Y=1041340
X4012 1973 1969 1 1973 1969 1987 2 MOAI1S $T=319920 971160 0 0 $X=319920 $Y=970780
X4013 1985 1986 1 1977 2001 2003 2 MOAI1S $T=323020 940920 1 0 $X=323020 $Y=935500
X4014 1984 1995 1 1984 1995 2017 2 MOAI1S $T=323640 1031640 0 0 $X=323640 $Y=1031260
X4015 1936 1915 1 1936 1915 2012 2 MOAI1S $T=323640 1051800 1 0 $X=323640 $Y=1046380
X4016 1939 1999 1 1939 2011 1990 2 MOAI1S $T=324260 1021560 1 0 $X=324260 $Y=1016140
X4017 2001 2002 1 1980 1985 2018 2 MOAI1S $T=324880 930840 1 0 $X=324880 $Y=925420
X4018 2000 2003 1 2000 2003 2033 2 MOAI1S $T=324880 951000 1 0 $X=324880 $Y=945580
X4019 121 130 1 121 2019 125 2 MOAI1S $T=331080 1082040 1 180 $X=327360 $Y=1081660
X4020 2002 2001 1 2018 2042 2060 2 MOAI1S $T=328600 930840 1 0 $X=328600 $Y=925420
X4021 1935 2044 1 1935 2058 2070 2 MOAI1S $T=330460 1021560 1 0 $X=330460 $Y=1016140
X4022 2035 2026 1 2035 2026 2058 2 MOAI1S $T=330460 1061880 0 0 $X=330460 $Y=1061500
X4023 2038 2018 1 2038 2018 2083 2 MOAI1S $T=333560 930840 0 0 $X=333560 $Y=930460
X4024 2040 2082 1 2040 2082 2101 2 MOAI1S $T=336040 910680 1 0 $X=336040 $Y=905260
X4025 2071 1906 1 2020 70 2086 2 MOAI1S $T=340380 940920 1 180 $X=336660 $Y=940540
X4026 2041 2095 1 2041 2095 2144 2 MOAI1S $T=339760 910680 0 0 $X=339760 $Y=910300
X4027 2111 2110 1 2111 2104 2140 2 MOAI1S $T=342240 1071960 1 0 $X=342240 $Y=1066540
X4028 2136 1982 1 2136 1982 2158 2 MOAI1S $T=343480 981240 1 0 $X=343480 $Y=975820
X4029 2151 2156 1 2151 2108 2145 2 MOAI1S $T=348440 1051800 1 180 $X=344720 $Y=1051420
X4030 2153 2059 1 2153 2059 2152 2 MOAI1S $T=349680 951000 0 180 $X=345960 $Y=945580
X4031 2157 2154 1 2157 2154 2133 2 MOAI1S $T=350300 961080 0 180 $X=346580 $Y=955660
X4032 2121 2163 1 2121 2163 2178 2 MOAI1S $T=347820 1041720 0 0 $X=347820 $Y=1041340
X4033 2151 2179 1 2151 2155 2164 2 MOAI1S $T=352160 1051800 0 180 $X=348440 $Y=1046380
X4034 2149 2167 1 2149 2183 2180 2 MOAI1S $T=349060 1021560 1 0 $X=349060 $Y=1016140
X4035 2200 2188 1 2176 2059 2073 2 MOAI1S $T=353400 951000 0 180 $X=349680 $Y=945580
X4036 2149 2190 1 2149 2203 2208 2 MOAI1S $T=351540 1041720 0 0 $X=351540 $Y=1041340
X4037 2199 2205 1 2199 2205 2234 2 MOAI1S $T=354020 920760 1 0 $X=354020 $Y=915340
X4038 173 2170 1 173 2170 2205 2 MOAI1S $T=359600 910680 0 180 $X=355880 $Y=905260
X4039 1926 2220 1 1926 2220 2239 2 MOAI1S $T=355880 1051800 1 0 $X=355880 $Y=1046380
X4040 2210 2016 1 2210 2016 2218 2 MOAI1S $T=360220 1021560 0 180 $X=356500 $Y=1016140
X4041 2240 2075 1 2240 2075 2247 2 MOAI1S $T=360220 961080 1 0 $X=360220 $Y=955660
X4042 2151 2264 1 2151 2251 2227 2 MOAI1S $T=366420 1051800 1 180 $X=362700 $Y=1051420
X4043 105 166 1 2248 172 2265 2 MOAI1S $T=369520 940920 0 180 $X=365800 $Y=935500
X4044 2276 2271 1 2276 2271 2249 2 MOAI1S $T=369520 951000 1 180 $X=365800 $Y=950620
X4045 2229 2262 1 2263 2075 2309 2 MOAI1S $T=365800 961080 1 0 $X=365800 $Y=955660
X4046 2322 2318 1 2322 2318 2314 2 MOAI1S $T=375720 940920 0 180 $X=372000 $Y=935500
X4047 2327 2323 1 2327 2323 2320 2 MOAI1S $T=376340 951000 0 180 $X=372620 $Y=945580
X4048 105 196 1 2248 188 2351 2 MOAI1S $T=381920 920760 1 180 $X=378200 $Y=920380
X4049 2371 2316 1 2371 2316 2395 2 MOAI1S $T=381300 940920 1 0 $X=381300 $Y=935500
X4050 116 196 1 201 203 2400 2 MOAI1S $T=383780 910680 0 0 $X=383780 $Y=910300
X4051 2417 2234 1 2417 2234 2429 2 MOAI1S $T=388120 910680 0 0 $X=388120 $Y=910300
X4052 2429 212 1 2429 212 216 2 MOAI1S $T=390600 900600 0 0 $X=390600 $Y=900220
X4053 2450 2459 1 2450 2445 2422 2 MOAI1S $T=394940 991320 0 180 $X=391220 $Y=985900
X4054 2398 2409 1 2398 2445 2423 2 MOAI1S $T=394940 1001400 1 180 $X=391220 $Y=1001020
X4055 2465 2474 1 2465 2445 2453 2 MOAI1S $T=398040 1021560 0 180 $X=394320 $Y=1016140
X4056 2463 2448 1 2463 2448 2471 2 MOAI1S $T=394940 940920 0 0 $X=394940 $Y=940540
X4057 2489 2117 1 2489 2117 2487 2 MOAI1S $T=402380 940920 1 180 $X=398660 $Y=940540
X4058 2515 2533 1 2515 2513 2508 2 MOAI1S $T=407340 991320 1 180 $X=403620 $Y=990940
X4059 2450 2324 1 2450 2513 2481 2 MOAI1S $T=408580 981240 0 180 $X=404860 $Y=975820
X4060 2564 2480 1 2564 2445 2543 2 MOAI1S $T=414160 961080 1 180 $X=410440 $Y=960700
X4061 2517 2585 1 2517 2601 2622 2 MOAI1S $T=414160 1001400 0 0 $X=414160 $Y=1001020
X4062 2486 2586 1 2486 2601 2599 2 MOAI1S $T=414160 1021560 1 0 $X=414160 $Y=1016140
X4063 2595 2605 1 2595 2445 2565 2 MOAI1S $T=418500 961080 1 180 $X=414780 $Y=960700
X4064 2607 2573 1 2607 2445 2594 2 MOAI1S $T=420360 971160 1 180 $X=416640 $Y=970780
X4065 2517 2606 1 2517 2513 2617 2 MOAI1S $T=416640 1001400 1 0 $X=416640 $Y=995980
X4066 2607 2499 1 2607 2513 2633 2 MOAI1S $T=417880 981240 1 0 $X=417880 $Y=975820
X4067 2564 2613 1 2564 2513 2628 2 MOAI1S $T=418500 961080 1 0 $X=418500 $Y=955660
X4068 2619 2656 1 2619 2513 2603 2 MOAI1S $T=426560 1001400 0 180 $X=422840 $Y=995980
X4069 2619 2657 1 2619 2601 2641 2 MOAI1S $T=426560 1011480 0 180 $X=422840 $Y=1006060
X4070 2607 2688 1 2607 2679 2659 2 MOAI1S $T=432140 971160 1 180 $X=428420 $Y=970780
X4071 2675 2695 1 2517 2679 2648 2 MOAI1S $T=433380 1001400 0 180 $X=429660 $Y=995980
X4072 2595 2708 1 2595 2650 2720 2 MOAI1S $T=434000 961080 0 0 $X=434000 $Y=960700
X4073 2515 2408 1 2515 2679 2725 2 MOAI1S $T=435860 1001400 1 0 $X=435860 $Y=995980
X4074 2718 2666 1 2718 2601 2733 2 MOAI1S $T=435860 1011480 0 0 $X=435860 $Y=1011100
X4075 2730 2731 1 2730 2650 2690 2 MOAI1S $T=441440 940920 1 180 $X=437720 $Y=940540
X4076 2564 2727 1 2564 2679 2739 2 MOAI1S $T=437720 961080 1 0 $X=437720 $Y=955660
X4077 2450 2754 1 2450 2679 2697 2 MOAI1S $T=445160 981240 0 180 $X=441440 $Y=975820
X4078 2730 2437 1 2730 2747 2719 2 MOAI1S $T=445780 940920 1 180 $X=442060 $Y=940540
X4079 2595 2780 1 2595 2747 2732 2 MOAI1S $T=448260 951000 1 180 $X=444540 $Y=950620
X4080 2748 2781 1 2619 2679 2756 2 MOAI1S $T=448260 991320 1 180 $X=444540 $Y=990940
X4081 2782 2792 1 2782 2650 2773 2 MOAI1S $T=450120 940920 1 180 $X=446400 $Y=940540
X4082 2718 2829 1 2718 2818 2787 2 MOAI1S $T=456940 1031640 0 180 $X=453220 $Y=1026220
X4083 2813 2837 1 2813 2805 2814 2 MOAI1S $T=458800 971160 0 180 $X=455080 $Y=965740
X4084 2823 2827 1 2823 2805 2845 2 MOAI1S $T=455080 1001400 0 0 $X=455080 $Y=1001020
X4085 2711 2831 1 2711 2805 2844 2 MOAI1S $T=455700 991320 1 0 $X=455700 $Y=985900
X4086 2810 2848 1 2810 2650 2868 2 MOAI1S $T=458800 961080 1 0 $X=458800 $Y=955660
X4087 2782 2558 1 2782 2747 2858 2 MOAI1S $T=459420 940920 0 0 $X=459420 $Y=940540
X4088 2810 2820 1 2810 2747 2863 2 MOAI1S $T=459420 951000 1 0 $X=459420 $Y=945580
X4089 2748 2865 1 2748 2805 2850 2 MOAI1S $T=463760 991320 0 180 $X=460040 $Y=985900
X4090 2812 2857 1 2812 2818 2870 2 MOAI1S $T=460660 1031640 1 0 $X=460660 $Y=1026220
X4091 2851 2871 1 2851 2818 2847 2 MOAI1S $T=465000 1001400 1 180 $X=461280 $Y=1001020
X4092 2711 2890 1 2711 2818 2885 2 MOAI1S $T=469340 1001400 1 180 $X=465620 $Y=1001020
X4093 2782 2915 1 2782 2906 2883 2 MOAI1S $T=473680 940920 1 180 $X=469960 $Y=940540
X4094 2812 2467 1 2812 2906 2922 2 MOAI1S $T=471200 971160 1 0 $X=471200 $Y=965740
X4095 2838 2917 1 2838 2805 2935 2 MOAI1S $T=471820 981240 0 0 $X=471820 $Y=980860
X4096 2942 2938 1 2810 2906 2899 2 MOAI1S $T=478020 951000 1 180 $X=474300 $Y=950620
X4097 2748 2903 1 2748 2818 2910 2 MOAI1S $T=478640 991320 1 180 $X=474920 $Y=990940
X4098 310 2920 1 306 2898 2877 2 MOAI1S $T=479260 1071960 1 180 $X=475540 $Y=1071580
X4099 2813 2943 1 2813 2818 2960 2 MOAI1S $T=476780 1031640 1 0 $X=476780 $Y=1026220
X4100 310 2973 1 306 2957 2972 2 MOAI1S $T=486700 1071960 0 180 $X=482980 $Y=1066540
X4101 310 2999 1 306 316 2981 2 MOAI1S $T=487940 1071960 1 180 $X=484220 $Y=1071580
X4102 310 3002 1 3004 320 3024 2 MOAI1S $T=486700 1071960 1 0 $X=486700 $Y=1066540
X4103 3005 3016 1 3005 2997 2967 2 MOAI1S $T=491660 1031640 0 180 $X=487940 $Y=1026220
X4104 260 3043 1 325 297 3003 2 MOAI1S $T=496620 900600 1 180 $X=492900 $Y=900220
X4105 3037 3046 1 3037 2997 3032 2 MOAI1S $T=496620 1031640 0 180 $X=492900 $Y=1026220
X4106 310 3029 1 306 326 3033 2 MOAI1S $T=497860 1071960 1 180 $X=494140 $Y=1071580
X4107 3059 3057 1 3004 327 3047 2 MOAI1S $T=499100 1061880 0 180 $X=495380 $Y=1056460
X4108 3060 2618 1 3060 295 3058 2 MOAI1S $T=501580 920760 1 180 $X=497860 $Y=920380
X4109 332 2996 1 3004 3027 3063 2 MOAI1S $T=502820 1041720 0 180 $X=499100 $Y=1036300
X4110 3069 3045 1 3069 334 3084 2 MOAI1S $T=500960 961080 0 0 $X=500960 $Y=960700
X4111 3059 3083 1 3077 3030 3074 2 MOAI1S $T=504680 1021560 1 180 $X=500960 $Y=1021180
X4112 2942 3082 1 2942 334 3094 2 MOAI1S $T=502820 951000 1 0 $X=502820 $Y=945580
X4113 3059 3100 1 3077 3080 3087 2 MOAI1S $T=507780 1041720 1 180 $X=504060 $Y=1041340
X4114 3005 2217 1 3005 3113 3078 2 MOAI1S $T=505920 981240 0 0 $X=505920 $Y=980860
X4115 3037 3105 1 3037 2601 3131 2 MOAI1S $T=506540 1011480 0 0 $X=506540 $Y=1011100
X4116 3059 3091 1 3077 3118 3120 2 MOAI1S $T=506540 1031640 1 0 $X=506540 $Y=1026220
X4117 3101 3110 1 3101 297 3119 2 MOAI1S $T=507160 910680 1 0 $X=507160 $Y=905260
X4118 3146 2165 1 3132 3113 3111 2 MOAI1S $T=514600 961080 0 180 $X=510880 $Y=955660
X4119 3141 353 1 3005 3123 3102 2 MOAI1S $T=514600 981240 1 180 $X=510880 $Y=980860
X4120 3132 3142 1 3132 334 3107 2 MOAI1S $T=515840 940920 1 180 $X=512120 $Y=940540
X4121 3106 3145 1 3106 3123 3124 2 MOAI1S $T=515840 1001400 0 180 $X=512120 $Y=995980
X4122 3121 3137 1 3121 2997 3148 2 MOAI1S $T=512120 1031640 1 0 $X=512120 $Y=1026220
X4123 3101 355 1 3101 3123 3168 2 MOAI1S $T=515840 910680 1 0 $X=515840 $Y=905260
X4124 3132 3162 1 3132 295 3130 2 MOAI1S $T=519560 940920 1 180 $X=515840 $Y=940540
X4125 3106 3152 1 3106 2997 3191 2 MOAI1S $T=515840 1031640 1 0 $X=515840 $Y=1026220
X4126 3139 3154 1 3139 295 3170 2 MOAI1S $T=516460 930840 1 0 $X=516460 $Y=925420
X4127 3169 2444 1 3169 3175 3109 2 MOAI1S $T=523280 971160 1 180 $X=519560 $Y=970780
X4128 3114 362 1 3114 3113 3172 2 MOAI1S $T=523280 981240 1 180 $X=519560 $Y=980860
X4129 3139 3179 1 3139 363 3204 2 MOAI1S $T=520180 920760 0 0 $X=520180 $Y=920380
X4130 3141 2545 1 3141 3175 3108 2 MOAI1S $T=525140 971160 0 180 $X=521420 $Y=965740
X4131 3190 2295 1 3190 2906 3184 2 MOAI1S $T=525760 940920 1 180 $X=522040 $Y=940540
X4132 3169 3198 1 3114 3209 3181 2 MOAI1S $T=523280 981240 0 0 $X=523280 $Y=980860
X4133 3121 3200 1 3121 3123 3210 2 MOAI1S $T=523280 1011480 1 0 $X=523280 $Y=1006060
X4134 365 3211 1 365 363 3186 2 MOAI1S $T=528240 910680 0 180 $X=524520 $Y=905260
X4135 3190 2392 1 3190 3175 3196 2 MOAI1S $T=529480 940920 1 180 $X=525760 $Y=940540
X4136 3231 374 1 3231 3219 3202 2 MOAI1S $T=533200 1011480 0 180 $X=529480 $Y=1006060
X4137 3240 3243 1 3240 334 3267 2 MOAI1S $T=533200 971160 1 0 $X=533200 $Y=965740
X4138 3245 3254 1 3245 3219 3230 2 MOAI1S $T=536920 1011480 0 180 $X=533200 $Y=1006060
X4139 3141 3247 1 3141 3259 3264 2 MOAI1S $T=533820 991320 1 0 $X=533820 $Y=985900
X4140 365 3263 1 3101 388 3273 2 MOAI1S $T=536300 910680 1 0 $X=536300 $Y=905260
X4141 3222 3288 1 3222 3209 3251 2 MOAI1S $T=543120 951000 0 180 $X=539400 $Y=945580
X4142 332 3285 1 3077 3297 394 2 MOAI1S $T=540640 910680 1 0 $X=540640 $Y=905260
X4143 3146 3300 1 3146 3280 3274 2 MOAI1S $T=544360 940920 1 180 $X=540640 $Y=940540
X4144 3303 397 1 3303 3277 3252 2 MOAI1S $T=546220 1011480 1 180 $X=542500 $Y=1011100
X4145 3309 2241 1 3309 3277 3317 2 MOAI1S $T=544360 1031640 0 0 $X=544360 $Y=1031260
X4146 401 3327 1 401 3176 3256 2 MOAI1S $T=546840 910680 1 0 $X=546840 $Y=905260
X4147 3303 3332 1 3303 3176 3342 2 MOAI1S $T=547460 1021560 0 0 $X=547460 $Y=1021180
X4148 3345 411 1 3345 3277 3340 2 MOAI1S $T=553660 1031640 1 180 $X=549940 $Y=1031260
X4149 3353 2257 1 3353 3277 3350 2 MOAI1S $T=554900 1011480 1 180 $X=551180 $Y=1011100
X4150 3358 3362 1 3358 388 3380 2 MOAI1S $T=553660 910680 1 0 $X=553660 $Y=905260
X4151 3369 3383 1 3369 3277 3366 2 MOAI1S $T=558620 1001400 0 180 $X=554900 $Y=995980
X4152 3378 2250 1 3378 3277 3302 2 MOAI1S $T=559860 1011480 0 180 $X=556140 $Y=1006060
X4153 3353 3415 1 3353 3259 3376 2 MOAI1S $T=563580 1011480 0 180 $X=559860 $Y=1006060
X4154 3373 2698 1 3373 3420 3428 2 MOAI1S $T=560480 971160 1 0 $X=560480 $Y=965740
X4155 3409 3422 1 3409 3259 3394 2 MOAI1S $T=564820 1001400 0 180 $X=561100 $Y=995980
X4156 3409 427 1 3409 3399 3379 2 MOAI1S $T=564820 1031640 1 180 $X=561100 $Y=1031260
X4157 3343 3425 1 3343 3259 3452 2 MOAI1S $T=563580 981240 0 0 $X=563580 $Y=980860
X4158 3343 3432 1 3343 3420 3442 2 MOAI1S $T=564820 961080 1 0 $X=564820 $Y=955660
X4159 3231 432 1 3231 3399 3439 2 MOAI1S $T=564820 1041720 1 0 $X=564820 $Y=1036300
X4160 3414 2626 1 3414 3175 3457 2 MOAI1S $T=567300 940920 0 0 $X=567300 $Y=940540
X4161 3321 3460 1 3321 3420 3447 2 MOAI1S $T=572260 971160 0 180 $X=568540 $Y=965740
X4162 3321 439 1 3321 3464 3453 2 MOAI1S $T=569780 1001400 1 0 $X=569780 $Y=995980
X4163 3458 3472 1 3458 3464 3433 2 MOAI1S $T=574740 991320 0 180 $X=571020 $Y=985900
X4164 3368 3504 1 3368 3464 3465 2 MOAI1S $T=582800 961080 0 180 $X=579080 $Y=955660
X4165 3496 464 1 3496 3464 3469 2 MOAI1S $T=583420 1001400 0 180 $X=579700 $Y=995980
X4166 3496 457 1 3496 3420 3523 2 MOAI1S $T=580320 971160 1 0 $X=580320 $Y=965740
X4167 3368 3506 1 3368 3399 3530 2 MOAI1S $T=580940 1031640 1 0 $X=580940 $Y=1026220
X4168 3414 3501 1 3414 3280 3522 2 MOAI1S $T=581560 940920 0 0 $X=581560 $Y=940540
X4169 3440 463 1 3440 3259 3525 2 MOAI1S $T=581560 981240 0 0 $X=581560 $Y=980860
X4170 3440 3515 1 3440 3464 3545 2 MOAI1S $T=582800 991320 1 0 $X=582800 $Y=985900
X4171 3516 3526 1 3516 3399 3537 2 MOAI1S $T=584040 1041720 1 0 $X=584040 $Y=1036300
X4172 3369 3555 1 3369 3464 3542 2 MOAI1S $T=593340 1001400 0 180 $X=589620 $Y=995980
X4173 3558 3562 1 3558 3420 3574 2 MOAI1S $T=592720 971160 1 0 $X=592720 $Y=965740
X4174 3558 3565 1 3558 3259 3572 2 MOAI1S $T=593340 981240 0 0 $X=593340 $Y=980860
X4175 507 509 1 514 3666 3671 2 MOAI1S $T=611320 1082040 0 0 $X=611320 $Y=1081660
X4176 507 3625 1 514 3633 3681 2 MOAI1S $T=611940 1082040 1 0 $X=611940 $Y=1076620
X4177 3647 515 1 3647 3676 3598 2 MOAI1S $T=613180 1011480 1 0 $X=613180 $Y=1006060
X4178 3679 3693 1 3679 3676 3672 2 MOAI1S $T=618760 991320 0 180 $X=615040 $Y=985900
X4179 3702 3505 1 3702 3676 3642 2 MOAI1S $T=621240 961080 1 180 $X=617520 $Y=960700
X4180 3704 526 1 3704 3676 3615 2 MOAI1S $T=621240 1011480 0 180 $X=617520 $Y=1006060
X4181 3726 532 1 3726 3676 3635 2 MOAI1S $T=624960 951000 1 180 $X=621240 $Y=950620
X4182 3657 3734 1 3657 529 3714 2 MOAI1S $T=624960 961080 1 180 $X=621240 $Y=960700
X4183 3746 3590 1 3746 3676 3727 2 MOAI1S $T=631780 991320 0 180 $X=628060 $Y=985900
X4184 3726 542 1 3726 3786 3792 2 MOAI1S $T=631780 940920 0 0 $X=631780 $Y=940540
X4185 546 548 1 546 529 3787 2 MOAI1S $T=637980 951000 1 180 $X=634260 $Y=950620
X4186 3657 549 1 3795 3786 3760 2 MOAI1S $T=637980 961080 1 180 $X=634260 $Y=960700
X4187 3647 3789 1 3813 3815 3818 2 MOAI1S $T=638600 1011480 1 0 $X=638600 $Y=1006060
X4188 3812 3594 1 3726 3280 3810 2 MOAI1S $T=643560 951000 0 180 $X=639840 $Y=945580
X4189 3679 560 1 3679 3815 3784 2 MOAI1S $T=643560 991320 0 180 $X=639840 $Y=985900
X4190 3704 3831 1 3704 3815 3844 2 MOAI1S $T=642940 1011480 1 0 $X=642940 $Y=1006060
X4191 3830 561 1 3830 3834 3850 2 MOAI1S $T=643560 981240 1 0 $X=643560 $Y=975820
X4192 3746 562 1 3839 3815 3857 2 MOAI1S $T=643560 991320 0 0 $X=643560 $Y=990940
X4193 3795 3618 1 3795 3846 3816 2 MOAI1S $T=651000 961080 0 180 $X=647280 $Y=955660
X4194 3830 3866 1 3830 3846 3856 2 MOAI1S $T=652240 971160 1 180 $X=648520 $Y=970780
X4195 3858 3634 1 3679 3867 3853 2 MOAI1S $T=654100 1001400 0 180 $X=650380 $Y=995980
X4196 3860 3877 1 3704 3867 3842 2 MOAI1S $T=654100 1011480 0 180 $X=650380 $Y=1006060
X4197 574 3825 1 534 3872 3894 2 MOAI1S $T=652860 920760 0 0 $X=652860 $Y=920380
X4198 3891 3855 1 582 3878 3916 2 MOAI1S $T=655960 1071960 0 0 $X=655960 $Y=1071580
X4199 3813 589 1 3813 3867 3886 2 MOAI1S $T=662160 1011480 1 180 $X=658440 $Y=1011100
X4200 3839 594 1 3839 3927 3958 2 MOAI1S $T=662160 1001400 1 0 $X=662160 $Y=995980
X4201 3812 3942 1 3812 3867 3960 2 MOAI1S $T=663400 940920 0 0 $X=663400 $Y=940540
X4202 3860 3659 1 3860 3927 3963 2 MOAI1S $T=664020 1011480 1 0 $X=664020 $Y=1006060
X4203 3938 3952 1 3938 3927 3981 2 MOAI1S $T=664640 1011480 0 0 $X=664640 $Y=1011100
X4204 587 3906 1 598 3965 3959 2 MOAI1S $T=664640 1082040 1 0 $X=664640 $Y=1076620
X4205 3940 3926 1 3830 3867 3977 2 MOAI1S $T=665260 971160 0 0 $X=665260 $Y=970780
X4206 3858 3583 1 3858 3846 3998 2 MOAI1S $T=667120 1001400 1 0 $X=667120 $Y=995980
X4207 626 4048 1 582 4025 4030 2 MOAI1S $T=681380 920760 1 180 $X=677660 $Y=920380
X4208 633 635 1 627 4010 4072 2 MOAI1S $T=684480 1082040 0 0 $X=684480 $Y=1081660
X4209 643 4092 1 630 4113 4062 2 MOAI1S $T=688200 1071960 0 0 $X=688200 $Y=1071580
X4210 4088 4133 1 4088 4146 4143 2 MOAI1S $T=694400 961080 1 0 $X=694400 $Y=955660
X4211 4080 3876 1 4080 4146 4156 2 MOAI1S $T=695640 951000 1 0 $X=695640 $Y=945580
X4212 4141 3827 1 4141 4137 4165 2 MOAI1S $T=696260 1001400 0 0 $X=696260 $Y=1001020
X4213 4066 4177 1 4066 4146 4157 2 MOAI1S $T=702460 991320 0 180 $X=698740 $Y=985900
X4214 4086 652 1 4171 4137 4185 2 MOAI1S $T=698740 1011480 1 0 $X=698740 $Y=1006060
X4215 4151 4183 1 4151 3834 4130 2 MOAI1S $T=704320 971160 1 180 $X=700600 $Y=970780
X4216 4192 4199 1 4192 3834 4188 2 MOAI1S $T=706800 961080 0 180 $X=703080 $Y=955660
X4217 4192 4200 1 4192 529 4172 2 MOAI1S $T=706800 961080 1 180 $X=703080 $Y=960700
X4218 4080 4204 1 4080 4193 4162 2 MOAI1S $T=707420 940920 1 180 $X=703700 $Y=940540
X4219 4055 658 1 4055 4193 4208 2 MOAI1S $T=703700 991320 1 0 $X=703700 $Y=985900
X4220 4151 4205 1 4151 529 4212 2 MOAI1S $T=705560 971160 0 0 $X=705560 $Y=970780
X4221 4192 4228 1 4192 4193 4207 2 MOAI1S $T=712380 951000 1 180 $X=708660 $Y=950620
X4222 4231 657 1 4247 4184 4255 2 MOAI1S $T=712380 1082040 0 0 $X=712380 $Y=1081660
X4223 4141 668 1 4141 4250 4213 2 MOAI1S $T=717960 1011480 1 180 $X=714240 $Y=1011100
X4224 4231 4214 1 4247 4260 4269 2 MOAI1S $T=715480 1082040 1 0 $X=715480 $Y=1076620
X4225 4087 672 1 4087 4193 4254 2 MOAI1S $T=720440 951000 1 180 $X=716720 $Y=950620
X4226 4171 4265 1 4171 4250 4173 2 MOAI1S $T=718580 1001400 0 0 $X=718580 $Y=1001020
X4227 4066 4267 1 4291 4250 4303 2 MOAI1S $T=721680 991320 1 0 $X=721680 $Y=985900
X4228 633 683 1 627 684 4316 2 MOAI1S $T=722920 1082040 0 0 $X=722920 $Y=1081660
X4229 633 4321 1 627 4338 4350 2 MOAI1S $T=727260 1082040 0 0 $X=727260 $Y=1081660
X4230 4297 4342 1 4297 4340 4379 2 MOAI1S $T=729740 981240 1 0 $X=729740 $Y=975820
X4231 4353 4359 1 4353 4340 4372 2 MOAI1S $T=731600 991320 1 0 $X=731600 $Y=985900
X4232 3975 4325 1 3975 4368 4375 2 MOAI1S $T=732220 940920 0 0 $X=732220 $Y=940540
X4233 4297 699 1 4297 3834 4393 2 MOAI1S $T=734080 971160 1 0 $X=734080 $Y=965740
X4234 4357 4071 1 4171 4380 4399 2 MOAI1S $T=734700 1001400 1 0 $X=734700 $Y=995980
X4235 701 704 1 701 4380 4374 2 MOAI1S $T=739040 951000 0 180 $X=735320 $Y=945580
X4236 4307 4298 1 4307 4340 4385 2 MOAI1S $T=740900 991320 0 180 $X=737180 $Y=985900
X4237 4227 4400 1 701 4368 4411 2 MOAI1S $T=739040 951000 1 0 $X=739040 $Y=945580
X4238 4381 3595 1 4381 4380 4422 2 MOAI1S $T=740280 971160 1 0 $X=740280 $Y=965740
X4239 4307 4415 1 4307 4421 4431 2 MOAI1S $T=742140 1011480 1 0 $X=742140 $Y=1006060
X4240 4381 4354 1 4381 4340 4430 2 MOAI1S $T=743380 981240 0 0 $X=743380 $Y=980860
X4241 4461 4491 1 4461 4368 4475 2 MOAI1S $T=760740 940920 1 180 $X=757020 $Y=940540
X4242 4513 4500 1 4513 4444 4439 2 MOAI1S $T=765080 1051800 0 180 $X=761360 $Y=1046380
X4243 4523 738 1 4523 4520 4451 2 MOAI1S $T=766940 1031640 1 180 $X=763220 $Y=1031260
X4244 4518 4458 1 4518 4380 4468 2 MOAI1S $T=767560 940920 1 180 $X=763840 $Y=940540
X4245 4528 4489 1 4528 4520 4453 2 MOAI1S $T=768180 1031640 0 180 $X=764460 $Y=1026220
X4246 4532 4384 1 4532 4531 4470 2 MOAI1S $T=769420 1021560 1 180 $X=765700 $Y=1021180
X4247 748 4553 1 748 747 4494 2 MOAI1S $T=771280 900600 1 180 $X=767560 $Y=900220
X4248 4539 749 1 4539 4368 4503 2 MOAI1S $T=771280 940920 1 180 $X=767560 $Y=940540
X4249 4547 750 1 4547 4380 4536 2 MOAI1S $T=771900 940920 0 180 $X=768180 $Y=935500
X4250 4532 4566 1 4532 4578 4480 2 MOAI1S $T=770660 1011480 1 0 $X=770660 $Y=1006060
X4251 735 4582 1 735 752 4567 2 MOAI1S $T=775000 900600 1 180 $X=771280 $Y=900220
X4252 4523 4530 1 4523 4562 4552 2 MOAI1S $T=775000 1021560 0 180 $X=771280 $Y=1016140
X4253 4522 4584 1 4522 4444 4537 2 MOAI1S $T=775000 1041720 1 180 $X=771280 $Y=1041340
X4254 4593 4599 1 4593 4578 4615 2 MOAI1S $T=775000 1011480 1 0 $X=775000 $Y=1006060
X4255 4518 4603 1 4518 4146 4495 2 MOAI1S $T=780580 920760 1 180 $X=776860 $Y=920380
X4256 4547 4588 1 4547 4578 4596 2 MOAI1S $T=781200 940920 0 180 $X=777480 $Y=935500
X4257 4729 4587 1 4729 810 4744 2 MOAI1S $T=801040 940920 0 180 $X=797320 $Y=935500
X4258 4709 4730 1 4709 4520 4707 2 MOAI1S $T=802280 1041720 0 180 $X=798560 $Y=1036300
X4259 4775 4779 1 4775 4578 4770 2 MOAI1S $T=804760 1011480 0 180 $X=801040 $Y=1006060
X4260 4794 4787 1 4780 810 4774 2 MOAI1S $T=805380 940920 0 180 $X=801660 $Y=935500
X4261 4729 4791 1 4729 4578 4691 2 MOAI1S $T=806000 951000 1 180 $X=802280 $Y=950620
X4262 4775 4798 1 4775 4531 4721 2 MOAI1S $T=806620 1021560 1 180 $X=802900 $Y=1021180
X4263 4709 4804 1 4775 4444 4776 2 MOAI1S $T=807240 1041720 1 180 $X=803520 $Y=1041340
X4264 4794 4811 1 4794 4578 4704 2 MOAI1S $T=808480 940920 1 180 $X=804760 $Y=940540
X4265 4853 4865 1 4853 4531 4802 2 MOAI1S $T=815920 1021560 0 180 $X=812200 $Y=1016140
X4266 4780 833 1 4695 4854 4851 2 MOAI1S $T=816540 951000 0 180 $X=812820 $Y=945580
X4267 4853 843 1 4853 4520 4835 2 MOAI1S $T=820880 1031640 0 180 $X=817160 $Y=1026220
X4268 4780 4900 1 4780 842 4875 2 MOAI1S $T=822740 930840 1 180 $X=819020 $Y=930460
X4269 4872 4771 1 4872 4520 4920 2 MOAI1S $T=823360 1041720 1 0 $X=823360 $Y=1036300
X4270 4902 4701 1 4902 4854 4940 2 MOAI1S $T=833280 951000 0 180 $X=829560 $Y=945580
X4271 4923 860 1 4923 4444 4969 2 MOAI1S $T=831420 1041720 0 0 $X=831420 $Y=1041340
X4272 4884 4950 1 4884 4444 4970 2 MOAI1S $T=831420 1051800 0 0 $X=831420 $Y=1051420
X4273 4902 4954 1 4902 4966 4963 2 MOAI1S $T=832040 940920 1 0 $X=832040 $Y=935500
X4274 4872 4957 1 4872 4531 4965 2 MOAI1S $T=832040 1021560 0 0 $X=832040 $Y=1021180
X4275 4977 5030 1 4977 4982 5002 2 MOAI1S $T=846300 1041720 0 180 $X=842580 $Y=1036300
X4276 5032 5115 1 5032 4968 5012 2 MOAI1S $T=861180 1021560 1 180 $X=857460 $Y=1021180
X4277 5007 5118 1 5007 4968 5111 2 MOAI1S $T=859940 1011480 0 0 $X=859940 $Y=1011100
X4278 5095 5119 1 5095 4982 5134 2 MOAI1S $T=859940 1041720 1 0 $X=859940 $Y=1036300
X4279 5095 903 1 5032 4531 5090 2 MOAI1S $T=867380 1021560 1 180 $X=863660 $Y=1021180
X4280 5149 5156 1 5149 4982 5096 2 MOAI1S $T=868000 1041720 0 180 $X=864280 $Y=1036300
X4281 5007 4978 1 5007 5173 5195 2 MOAI1S $T=869860 1021560 0 0 $X=869860 $Y=1021180
X4282 5213 5226 1 5213 5223 5167 2 MOAI1S $T=879780 1021560 1 180 $X=876060 $Y=1021180
X4283 5213 5234 1 5213 4982 5186 2 MOAI1S $T=880400 1041720 0 180 $X=876680 $Y=1036300
X4284 5138 5295 1 5138 929 5256 2 MOAI1S $T=889080 951000 1 180 $X=885360 $Y=950620
X4285 5245 930 1 5245 4982 5316 2 MOAI1S $T=885360 1041720 1 0 $X=885360 $Y=1036300
X4286 5275 5285 1 5275 5223 5312 2 MOAI1S $T=885980 1021560 0 0 $X=885980 $Y=1021180
X4287 5255 934 1 5255 4854 5286 2 MOAI1S $T=890940 940920 1 180 $X=887220 $Y=940540
X4288 5300 5307 1 5300 5173 5288 2 MOAI1S $T=890940 1031640 1 180 $X=887220 $Y=1031260
X4289 5296 5301 1 5296 5223 5252 2 MOAI1S $T=887840 1011480 1 0 $X=887840 $Y=1006060
X4290 5109 935 1 5109 929 5293 2 MOAI1S $T=892180 971160 1 180 $X=888460 $Y=970780
X4291 5284 5323 1 5284 5173 5332 2 MOAI1S $T=891560 1001400 1 0 $X=891560 $Y=995980
X4292 5296 5334 1 5296 5173 5346 2 MOAI1S $T=893420 1011480 1 0 $X=893420 $Y=1006060
X4293 5275 5347 1 5275 5173 5336 2 MOAI1S $T=897760 1021560 1 180 $X=894040 $Y=1021180
X4294 5263 943 1 5263 5173 5358 2 MOAI1S $T=895280 1001400 1 0 $X=895280 $Y=995980
X4295 5277 944 1 5277 4854 5361 2 MOAI1S $T=896520 951000 1 0 $X=896520 $Y=945580
X4296 5353 5376 1 5353 4968 5385 2 MOAI1S $T=900860 1011480 0 0 $X=900860 $Y=1011100
X4297 5277 952 1 5277 958 5394 2 MOAI1S $T=901480 940920 1 0 $X=901480 $Y=935500
X4298 5277 959 1 5277 4966 5368 2 MOAI1S $T=905200 940920 1 180 $X=901480 $Y=940540
X4299 5372 5384 1 5372 4968 5365 2 MOAI1S $T=905200 991320 1 180 $X=901480 $Y=990940
X4300 5275 953 1 5275 4968 5386 2 MOAI1S $T=901480 1021560 1 0 $X=901480 $Y=1016140
X4301 5372 5396 1 5372 5223 5355 2 MOAI1S $T=907680 971160 0 180 $X=903960 $Y=965740
X4302 5300 963 1 5300 4968 5421 2 MOAI1S $T=906440 1031640 0 0 $X=906440 $Y=1031260
X4303 5415 5392 1 5415 5223 5431 2 MOAI1S $T=912020 971160 1 0 $X=912020 $Y=965740
X4304 5255 5425 1 5255 4966 5438 2 MOAI1S $T=913880 951000 1 0 $X=913880 $Y=945580
X4305 5263 5426 1 5263 4966 5437 2 MOAI1S $T=913880 991320 0 0 $X=913880 $Y=990940
X4306 5415 5408 1 5415 4854 5462 2 MOAI1S $T=915740 971160 0 0 $X=915740 $Y=970780
X4307 5284 979 1 5284 4966 5439 2 MOAI1S $T=921320 991320 1 180 $X=917600 $Y=990940
X4308 5490 5476 1 5490 5486 5436 2 MOAI1S $T=927520 961080 1 180 $X=923800 $Y=960700
X4309 5523 5538 1 5523 5528 5502 2 MOAI1S $T=935580 991320 0 180 $X=931860 $Y=985900
X4310 5508 1013 1 5508 5528 5517 2 MOAI1S $T=939300 981240 1 180 $X=935580 $Y=980860
X4311 5527 5565 1 5527 5528 5600 2 MOAI1S $T=939920 981240 0 0 $X=939920 $Y=980860
X4312 5562 5607 1 5562 5528 5578 2 MOAI1S $T=946740 991320 0 180 $X=943020 $Y=985900
X4313 5678 5688 1 5678 5528 5673 2 MOAI1S $T=959760 991320 0 180 $X=956040 $Y=985900
X4314 1029 5716 1 1029 1045 5703 2 MOAI1S $T=964720 910680 0 180 $X=961000 $Y=905260
X4315 5721 5587 1 5721 5757 5737 2 MOAI1S $T=968440 1001400 1 0 $X=968440 $Y=995980
X4316 5779 5775 1 5779 5757 5802 2 MOAI1S $T=977740 991320 0 0 $X=977740 $Y=990940
X4317 5796 5674 1 5796 5757 5807 2 MOAI1S $T=980840 1001400 0 0 $X=980840 $Y=1001020
X4318 5828 1074 1 5810 958 5793 2 MOAI1S $T=987040 940920 1 180 $X=983320 $Y=940540
X4319 5829 5837 1 5829 5757 5814 2 MOAI1S $T=992000 1011480 0 180 $X=988280 $Y=1006060
X4320 5810 5846 1 5810 929 5825 2 MOAI1S $T=993240 971160 1 180 $X=989520 $Y=970780
X4321 5810 1083 1 5810 5486 5789 2 MOAI1S $T=993860 961080 0 180 $X=990140 $Y=955660
X4322 5856 5861 1 5856 5852 5838 2 MOAI1S $T=996340 940920 1 180 $X=992620 $Y=940540
X4323 5857 5830 1 5857 5757 5815 2 MOAI1S $T=996340 1011480 0 180 $X=992620 $Y=1006060
X4324 5858 5869 1 5858 929 5848 2 MOAI1S $T=998200 971160 1 180 $X=994480 $Y=970780
X4325 1077 5871 1 1077 1087 5831 2 MOAI1S $T=999440 900600 1 180 $X=995720 $Y=900220
X4326 5856 5873 1 5856 5486 5850 2 MOAI1S $T=999440 961080 0 180 $X=995720 $Y=955660
X4327 5829 5875 1 5829 5866 5834 2 MOAI1S $T=999440 981240 1 180 $X=995720 $Y=980860
X4328 5857 5876 1 5857 5866 5844 2 MOAI1S $T=999440 991320 1 180 $X=995720 $Y=990940
X4329 5897 5909 1 5897 5757 5880 2 MOAI1S $T=1004400 1011480 0 180 $X=1000680 $Y=1006060
X4330 5905 1102 1 5905 5852 5817 2 MOAI1S $T=1005640 930840 1 180 $X=1001920 $Y=930460
X4331 5915 5931 1 5915 1099 5908 2 MOAI1S $T=1006880 971160 1 180 $X=1003160 $Y=970780
X4332 5897 1105 1 5897 5866 5935 2 MOAI1S $T=1004400 1001400 1 0 $X=1004400 $Y=995980
X4333 5918 5862 1 5918 1099 5912 2 MOAI1S $T=1008740 981240 0 180 $X=1005020 $Y=975820
X4334 5921 5835 1 5921 1109 5878 2 MOAI1S $T=1009360 920760 0 180 $X=1005640 $Y=915340
X4335 5915 5949 1 5915 1109 5914 2 MOAI1S $T=1010600 940920 1 180 $X=1006880 $Y=940540
X4336 5930 5946 1 5930 958 5954 2 MOAI1S $T=1007500 930840 0 0 $X=1007500 $Y=930460
X4337 5930 1117 1 5930 5486 5926 2 MOAI1S $T=1011220 961080 0 180 $X=1007500 $Y=955660
X4338 1077 1119 1 1077 1109 5966 2 MOAI1S $T=1009980 910680 0 0 $X=1009980 $Y=910300
X4339 5921 5988 1 5921 1127 5967 2 MOAI1S $T=1016800 920760 0 180 $X=1013080 $Y=915340
X4340 5986 5997 1 5986 5983 5970 2 MOAI1S $T=1018040 1011480 0 180 $X=1014320 $Y=1006060
X4341 6000 1136 1 6000 5852 5981 2 MOAI1S $T=1019900 940920 0 180 $X=1016180 $Y=935500
X4342 6027 1147 1 6027 5866 6021 2 MOAI1S $T=1025480 991320 1 180 $X=1021760 $Y=990940
X4343 6026 5992 1 6026 6039 6048 2 MOAI1S $T=1022380 961080 1 0 $X=1022380 $Y=955660
X4344 6026 6033 1 6026 1099 6042 2 MOAI1S $T=1023000 981240 1 0 $X=1023000 $Y=975820
X4345 1146 6038 1 1146 1127 6056 2 MOAI1S $T=1024240 910680 0 0 $X=1024240 $Y=910300
X4346 6027 6057 1 6027 5983 6043 2 MOAI1S $T=1029820 1011480 0 180 $X=1026100 $Y=1006060
X4347 6045 6058 1 6045 6039 6067 2 MOAI1S $T=1028580 961080 1 0 $X=1028580 $Y=955660
X4348 1154 6070 1 1154 1127 6053 2 MOAI1S $T=1032920 910680 1 180 $X=1029200 $Y=910300
X4349 6045 1153 1 6045 6071 6077 2 MOAI1S $T=1029200 940920 0 0 $X=1029200 $Y=940540
X4350 6063 6072 1 6063 6060 6047 2 MOAI1S $T=1032920 981240 1 180 $X=1029200 $Y=980860
X4351 6081 1159 1 6081 6071 6084 2 MOAI1S $T=1037880 951000 0 180 $X=1034160 $Y=945580
X4352 6080 6089 1 6080 5983 6106 2 MOAI1S $T=1034160 1001400 0 0 $X=1034160 $Y=1001020
X4353 6088 6044 1 6088 5866 6103 2 MOAI1S $T=1034780 930840 0 0 $X=1034780 $Y=930460
X4354 6091 6112 1 6091 6101 6087 2 MOAI1S $T=1039740 971160 0 180 $X=1036020 $Y=965740
X4355 6091 6030 1 6091 6060 6085 2 MOAI1S $T=1039740 981240 1 180 $X=1036020 $Y=980860
X4356 6116 6123 1 6116 5983 6104 2 MOAI1S $T=1042220 1011480 1 180 $X=1038500 $Y=1011100
X4357 6119 6100 1 6119 6071 6107 2 MOAI1S $T=1044700 951000 0 180 $X=1040980 $Y=945580
X4358 6145 6140 1 6125 5866 6121 2 MOAI1S $T=1045940 940920 0 180 $X=1042220 $Y=935500
X4359 6158 1179 1 6158 5983 6166 2 MOAI1S $T=1047180 1011480 0 0 $X=1047180 $Y=1011100
X4360 6142 1181 1 6142 6101 6094 2 MOAI1S $T=1048420 971160 0 0 $X=1048420 $Y=970780
X4361 6142 6170 1 6142 6060 6184 2 MOAI1S $T=1050900 991320 1 0 $X=1050900 $Y=985900
X4362 1188 1190 1 1188 6071 6177 2 MOAI1S $T=1056480 900600 1 180 $X=1052760 $Y=900220
X4363 6145 6214 1 6145 6206 6198 2 MOAI1S $T=1062060 940920 1 180 $X=1058340 $Y=940540
X4364 6190 6157 1 6190 6206 6217 2 MOAI1S $T=1058960 961080 0 0 $X=1058960 $Y=960700
X4365 6201 6219 1 6201 6101 6207 2 MOAI1S $T=1062680 971160 1 180 $X=1058960 $Y=970780
X4366 6197 1197 1 6197 6206 6229 2 MOAI1S $T=1059580 930840 1 0 $X=1059580 $Y=925420
X4367 6186 6235 1 6186 6206 6252 2 MOAI1S $T=1062680 930840 0 0 $X=1062680 $Y=930460
X4368 6181 1209 1 6181 6206 6245 2 MOAI1S $T=1070120 961080 0 180 $X=1066400 $Y=955660
X4369 6202 6262 1 6202 6101 6278 2 MOAI1S $T=1067020 971160 0 0 $X=1067020 $Y=970780
X4370 6168 6275 1 6168 6206 6286 2 MOAI1S $T=1070120 940920 1 0 $X=1070120 $Y=935500
X4371 1210 6285 1 1210 6071 6268 2 MOAI1S $T=1075080 910680 0 180 $X=1071360 $Y=905260
X4372 6202 6289 1 6202 6299 6301 2 MOAI1S $T=1074460 981240 0 0 $X=1074460 $Y=980860
X4373 6255 6306 1 6255 6299 6318 2 MOAI1S $T=1078180 981240 1 0 $X=1078180 $Y=975820
X4374 6303 1223 1 6303 6316 6258 2 MOAI1S $T=1078180 991320 0 0 $X=1078180 $Y=990940
X4375 6181 6308 1 6181 6299 6326 2 MOAI1S $T=1078800 961080 1 0 $X=1078800 $Y=955660
X4376 6190 1224 1 6190 6299 6327 2 MOAI1S $T=1078800 971160 1 0 $X=1078800 $Y=965740
X4377 6145 1228 1 6145 6315 6307 2 MOAI1S $T=1083760 940920 1 180 $X=1080040 $Y=940540
X4378 6290 1227 1 6290 6316 6270 2 MOAI1S $T=1080660 1001400 0 0 $X=1080660 $Y=1001020
X4379 6197 6334 1 6197 6315 6296 2 MOAI1S $T=1086240 930840 0 180 $X=1082520 $Y=925420
X4380 6290 6335 1 6290 6060 6314 2 MOAI1S $T=1086240 981240 0 180 $X=1082520 $Y=975820
X4381 6168 6361 1 6168 6315 6374 2 MOAI1S $T=1089340 940920 0 0 $X=1089340 $Y=940540
X4382 6186 6341 1 6186 6315 6377 2 MOAI1S $T=1089960 930840 1 0 $X=1089960 $Y=925420
X4383 6370 6375 1 6370 6316 6319 2 MOAI1S $T=1093680 1001400 1 180 $X=1089960 $Y=1001020
X4384 6303 6393 1 6303 6060 6356 2 MOAI1S $T=1096780 981240 1 180 $X=1093060 $Y=980860
X4385 6359 6384 1 6359 6399 6372 2 MOAI1S $T=1093680 991320 0 0 $X=1093680 $Y=990940
X4386 6415 6420 1 6415 6399 6410 2 MOAI1S $T=1101740 1001400 1 180 $X=1098020 $Y=1001020
X4387 6415 1258 1 6415 6426 6429 2 MOAI1S $T=1099880 971160 0 0 $X=1099880 $Y=970780
X4388 6370 1263 1 6370 6426 6404 2 MOAI1S $T=1104840 981240 0 180 $X=1101120 $Y=975820
X4389 6359 6449 1 6359 6426 6481 2 MOAI1S $T=1108560 981240 1 0 $X=1108560 $Y=975820
X4390 6408 6467 1 6408 6426 6496 2 MOAI1S $T=1109180 971160 1 0 $X=1109180 $Y=965740
X4391 6408 6479 1 6408 6468 6462 2 MOAI1S $T=1112900 1001400 0 180 $X=1109180 $Y=995980
X4392 6255 6490 1 6255 6426 6507 2 MOAI1S $T=1112900 981240 1 0 $X=1112900 $Y=975820
X4393 6486 6519 1 6486 6468 6523 2 MOAI1S $T=1120960 991320 0 0 $X=1120960 $Y=990940
X4394 6510 6526 1 6510 6426 6531 2 MOAI1S $T=1124680 971160 0 0 $X=1124680 $Y=970780
X4395 6510 6522 1 6510 6468 6529 2 MOAI1S $T=1125300 991320 0 0 $X=1125300 $Y=990940
X4396 1474 2 1428 23 1 NR2 $T=246140 920760 1 0 $X=246140 $Y=915340
X4397 1507 2 1489 1545 1 NR2 $T=254820 940920 1 0 $X=254820 $Y=935500
X4398 1567 2 1555 1534 1 NR2 $T=259780 1041720 0 180 $X=257920 $Y=1036300
X4399 39 2 1483 1560 1 NR2 $T=261640 1021560 0 180 $X=259780 $Y=1016140
X4400 1555 2 1585 1579 1 NR2 $T=259780 1051800 1 0 $X=259780 $Y=1046380
X4401 1601 2 1597 1570 1 NR2 $T=263500 961080 0 180 $X=261640 $Y=955660
X4402 1520 2 1494 1646 1 NR2 $T=262260 940920 1 0 $X=262260 $Y=935500
X4403 1612 2 1572 1591 1 NR2 $T=265360 1021560 1 180 $X=263500 $Y=1021180
X4404 1613 2 1605 1602 1 NR2 $T=266600 1041720 1 180 $X=264740 $Y=1041340
X4405 1597 2 1623 1610 1 NR2 $T=265360 961080 1 0 $X=265360 $Y=955660
X4406 47 2 1589 38 1 NR2 $T=268460 930840 0 180 $X=266600 $Y=925420
X4407 49 2 1596 47 1 NR2 $T=268460 940920 1 180 $X=266600 $Y=940540
X4408 48 2 44 47 1 NR2 $T=267220 910680 1 0 $X=267220 $Y=905260
X4409 50 2 1604 55 1 NR2 $T=269080 920760 1 0 $X=269080 $Y=915340
X4410 39 2 1584 1643 1 NR2 $T=269080 1021560 1 0 $X=269080 $Y=1016140
X4411 51 2 1524 1643 1 NR2 $T=272180 1021560 1 180 $X=270320 $Y=1021180
X4412 51 2 1640 1657 1 NR2 $T=270320 1031640 1 0 $X=270320 $Y=1026220
X4413 48 2 1654 57 1 NR2 $T=274040 920760 1 0 $X=274040 $Y=915340
X4414 1669 2 1580 1676 1 NR2 $T=274040 1051800 0 0 $X=274040 $Y=1051420
X4415 1653 2 1682 1658 1 NR2 $T=278380 1082040 1 180 $X=276520 $Y=1081660
X4416 57 2 1703 59 1 NR2 $T=279620 910680 0 180 $X=277760 $Y=905260
X4417 1696 2 1698 1700 1 NR2 $T=277760 971160 1 0 $X=277760 $Y=965740
X4418 49 2 1702 57 1 NR2 $T=279620 940920 0 0 $X=279620 $Y=940540
X4419 57 2 1662 38 1 NR2 $T=280860 940920 1 0 $X=280860 $Y=935500
X4420 1737 2 1694 55 1 NR2 $T=283340 910680 1 180 $X=281480 $Y=910300
X4421 57 2 1738 1737 1 NR2 $T=281480 920760 0 0 $X=281480 $Y=920380
X4422 39 2 1733 1657 1 NR2 $T=283340 1021560 1 0 $X=283340 $Y=1016140
X4423 1718 2 1720 1726 1 NR2 $T=285200 1051800 0 180 $X=283340 $Y=1046380
X4424 49 2 1727 1746 1 NR2 $T=284580 961080 0 0 $X=284580 $Y=960700
X4425 1758 2 1718 1671 1 NR2 $T=287060 1051800 0 180 $X=285200 $Y=1046380
X4426 1746 2 1750 1737 1 NR2 $T=288300 930840 1 180 $X=286440 $Y=930460
X4427 1737 2 1744 63 1 NR2 $T=286440 940920 1 0 $X=286440 $Y=935500
X4428 1746 2 1747 1734 1 NR2 $T=288920 961080 1 180 $X=287060 $Y=960700
X4429 1746 2 1457 73 1 NR2 $T=288300 910680 0 0 $X=288300 $Y=910300
X4430 1762 2 1520 1771 1 NR2 $T=288920 930840 0 0 $X=288920 $Y=930460
X4431 1778 2 1715 63 1 NR2 $T=290780 961080 0 180 $X=288920 $Y=955660
X4432 1772 2 1633 1790 1 NR2 $T=290160 961080 0 0 $X=290160 $Y=960700
X4433 1784 2 1735 1757 1 NR2 $T=292020 951000 0 0 $X=292020 $Y=950620
X4434 1612 2 1779 1657 1 NR2 $T=292020 1021560 0 0 $X=292020 $Y=1021180
X4435 66 2 1729 63 1 NR2 $T=293260 920760 1 0 $X=293260 $Y=915340
X4436 1813 2 1795 63 1 NR2 $T=295740 930840 0 180 $X=293880 $Y=925420
X4437 1746 2 1805 1813 1 NR2 $T=295120 920760 1 0 $X=295120 $Y=915340
X4438 69 2 1725 70 1 NR2 $T=297600 910680 1 0 $X=297600 $Y=905260
X4439 70 2 1798 71 1 NR2 $T=297600 930840 1 0 $X=297600 $Y=925420
X4440 73 2 1840 63 1 NR2 $T=300080 920760 0 180 $X=298220 $Y=915340
X4441 1831 2 1848 1847 1 NR2 $T=298220 1051800 1 0 $X=298220 $Y=1046380
X4442 1849 2 1801 1850 1 NR2 $T=299460 1061880 0 0 $X=299460 $Y=1061500
X4443 1853 2 1789 1818 1 NR2 $T=300080 930840 0 0 $X=300080 $Y=930460
X4444 1772 2 1786 71 1 NR2 $T=300700 961080 1 0 $X=300700 $Y=955660
X4445 1868 2 1860 1790 1 NR2 $T=302560 961080 1 180 $X=300700 $Y=960700
X4446 1869 2 1855 1831 1 NR2 $T=303800 1041720 0 180 $X=301940 $Y=1036300
X4447 77 2 1864 1887 1 NR2 $T=302560 910680 1 0 $X=302560 $Y=905260
X4448 70 2 1748 1871 1 NR2 $T=302560 920760 1 0 $X=302560 $Y=915340
X4449 77 2 1803 81 1 NR2 $T=302560 920760 0 0 $X=302560 $Y=920380
X4450 1874 2 1875 63 1 NR2 $T=304420 961080 0 180 $X=302560 $Y=955660
X4451 1862 2 1884 1829 1 NR2 $T=302560 981240 1 0 $X=302560 $Y=975820
X4452 1612 2 1879 1863 1 NR2 $T=304420 1031640 1 180 $X=302560 $Y=1031260
X4453 1869 2 1899 1848 1 NR2 $T=304420 1041720 1 180 $X=302560 $Y=1041340
X4454 1790 2 1842 1880 1 NR2 $T=303180 951000 0 0 $X=303180 $Y=950620
X4455 1868 2 1819 1871 1 NR2 $T=303180 961080 0 0 $X=303180 $Y=960700
X4456 1898 2 1869 1768 1 NR2 $T=305660 1041720 0 180 $X=303800 $Y=1036300
X4457 80 2 82 1887 1 NR2 $T=304420 900600 0 0 $X=304420 $Y=900220
X4458 80 2 1714 81 1 NR2 $T=306280 920760 0 180 $X=304420 $Y=915340
X4459 1880 2 1861 71 1 NR2 $T=304420 961080 1 0 $X=304420 $Y=955660
X4460 1911 2 1839 84 1 NR2 $T=308140 910680 0 180 $X=306280 $Y=905260
X4461 1880 2 1894 1871 1 NR2 $T=306280 951000 0 0 $X=306280 $Y=950620
X4462 1917 2 1811 71 1 NR2 $T=310000 961080 0 180 $X=308140 $Y=955660
X4463 1911 2 1909 1887 1 NR2 $T=309380 910680 1 0 $X=309380 $Y=905260
X4464 1911 2 86 97 1 NR2 $T=310000 900600 0 0 $X=310000 $Y=900220
X4465 1921 2 1876 1871 1 NR2 $T=311860 961080 1 180 $X=310000 $Y=960700
X4466 1821 2 1930 1914 1 NR2 $T=310000 1041720 0 0 $X=310000 $Y=1041340
X4467 102 2 1925 71 1 NR2 $T=313720 910680 0 180 $X=311860 $Y=905260
X4468 1930 2 1936 1901 1 NR2 $T=312480 1051800 1 0 $X=312480 $Y=1046380
X4469 97 2 1743 96 1 NR2 $T=316200 920760 0 180 $X=314340 $Y=915340
X4470 97 2 1942 99 1 NR2 $T=314960 910680 1 0 $X=314960 $Y=905260
X4471 96 2 1872 1887 1 NR2 $T=315580 920760 0 0 $X=315580 $Y=920380
X4472 99 2 1919 84 1 NR2 $T=316820 910680 1 0 $X=316820 $Y=905260
X4473 110 2 89 1887 1 NR2 $T=318680 910680 1 180 $X=316820 $Y=910300
X4474 1778 2 1959 1880 1 NR2 $T=316820 951000 0 0 $X=316820 $Y=950620
X4475 1778 2 1955 1868 1 NR2 $T=316820 961080 0 0 $X=316820 $Y=960700
X4476 113 2 1931 1868 1 NR2 $T=320540 961080 1 180 $X=318680 $Y=960700
X4477 1921 2 1986 1778 1 NR2 $T=321780 951000 0 180 $X=319920 $Y=945580
X4478 61 2 1975 1972 1 NR2 $T=321780 951000 1 180 $X=319920 $Y=950620
X4479 1921 2 1977 61 1 NR2 $T=320540 940920 1 0 $X=320540 $Y=935500
X4480 1974 2 1980 1917 1 NR2 $T=321160 930840 0 0 $X=321160 $Y=930460
X4481 1921 2 1973 1734 1 NR2 $T=321160 961080 0 0 $X=321160 $Y=960700
X4482 77 2 2001 1974 1 NR2 $T=322400 930840 1 0 $X=322400 $Y=925420
X4483 77 2 1985 61 1 NR2 $T=323020 930840 0 0 $X=323020 $Y=930460
X4484 61 2 2002 80 1 NR2 $T=325500 920760 1 180 $X=323640 $Y=920380
X4485 1772 2 1992 1734 1 NR2 $T=325500 971160 0 180 $X=323640 $Y=965740
X4486 1974 2 2006 110 1 NR2 $T=324260 920760 1 0 $X=324260 $Y=915340
X4487 61 2 1991 110 1 NR2 $T=326120 910680 1 0 $X=326120 $Y=905260
X4488 1974 2 2009 70 1 NR2 $T=326120 910680 0 0 $X=326120 $Y=910300
X4489 1772 2 2015 2020 1 NR2 $T=327360 961080 1 0 $X=327360 $Y=955660
X4490 1972 2 2022 1734 1 NR2 $T=329220 961080 1 180 $X=327360 $Y=960700
X4491 1917 2 2000 1734 1 NR2 $T=327980 930840 0 0 $X=327980 $Y=930460
X4492 1874 2 2028 1972 1 NR2 $T=331080 961080 0 180 $X=329220 $Y=955660
X4493 2020 2 2048 1972 1 NR2 $T=329220 971160 1 0 $X=329220 $Y=965740
X4494 1968 2 2038 1734 1 NR2 $T=332320 930840 1 180 $X=330460 $Y=930460
X4495 1921 2 2046 2020 1 NR2 $T=331080 951000 1 0 $X=331080 $Y=945580
X4496 1772 2 2061 1874 1 NR2 $T=331080 951000 0 0 $X=331080 $Y=950620
X4497 1921 2 2045 1874 1 NR2 $T=331080 961080 1 0 $X=331080 $Y=955660
X4498 2046 2 2047 2028 1 NR2 $T=332940 961080 1 180 $X=331080 $Y=960700
X4499 2054 2 2035 2021 1 NR2 $T=332940 1071960 0 180 $X=331080 $Y=1066540
X4500 2020 2 2065 1968 1 NR2 $T=334800 940920 0 180 $X=332940 $Y=935500
X4501 1874 2 2067 1868 1 NR2 $T=334800 961080 0 180 $X=332940 $Y=955660
X4502 2072 2 2062 2047 1 NR2 $T=334800 961080 1 180 $X=332940 $Y=960700
X4503 1874 2 2092 1917 1 NR2 $T=334800 951000 0 0 $X=334800 $Y=950620
X4504 2027 2 2021 2079 1 NR2 $T=334800 1071960 1 0 $X=334800 $Y=1066540
X4505 2020 2 2085 1917 1 NR2 $T=339140 951000 0 180 $X=337280 $Y=945580
X4506 2061 2 2105 2085 1 NR2 $T=338520 961080 1 0 $X=338520 $Y=955660
X4507 2112 2 2113 2076 1 NR2 $T=339760 930840 1 0 $X=339760 $Y=925420
X4508 2098 2 145 2134 1 NR2 $T=342240 1082040 1 0 $X=342240 $Y=1076620
X4509 2125 2 2132 2105 1 NR2 $T=344720 961080 0 180 $X=342860 $Y=955660
X4510 2121 2 2130 2129 1 NR2 $T=345340 1041720 1 0 $X=345340 $Y=1036300
X4511 160 2 2141 73 1 NR2 $T=349060 920760 1 180 $X=347200 $Y=920380
X4512 2136 2 2173 1982 1 NR2 $T=350920 981240 0 180 $X=349060 $Y=975820
X4513 2121 2 2174 2159 1 NR2 $T=349060 1021560 0 0 $X=349060 $Y=1021180
X4514 2174 2 2191 2161 1 NR2 $T=350920 1031640 0 180 $X=349060 $Y=1026220
X4515 113 2 2157 171 1 NR2 $T=352160 961080 1 0 $X=352160 $Y=955660
X4516 2177 2 2201 2204 1 NR2 $T=352160 1001400 0 0 $X=352160 $Y=1001020
X4517 2182 2 2197 2016 1 NR2 $T=352160 1021560 0 0 $X=352160 $Y=1021180
X4518 169 2 2188 2215 1 NR2 $T=354020 940920 0 0 $X=354020 $Y=940540
X4519 169 2 2143 172 1 NR2 $T=355260 940920 1 0 $X=355260 $Y=935500
X4520 1926 2 2211 2194 1 NR2 $T=355260 1041720 0 0 $X=355260 $Y=1041340
X4521 1790 2 2229 2215 1 NR2 $T=357740 940920 0 0 $X=357740 $Y=940540
X4522 1790 2 2223 171 1 NR2 $T=357740 961080 1 0 $X=357740 $Y=955660
X4523 2052 2 2252 73 1 NR2 $T=363320 920760 0 0 $X=363320 $Y=920380
X4524 2248 2 2228 2215 1 NR2 $T=363320 940920 1 0 $X=363320 $Y=935500
X4525 2248 2 2200 182 1 NR2 $T=363320 940920 0 0 $X=363320 $Y=940540
X4526 2248 2 2238 171 1 NR2 $T=363320 951000 1 0 $X=363320 $Y=945580
X4527 174 2 2253 172 1 NR2 $T=365180 940920 0 0 $X=365180 $Y=940540
X4528 81 2 2269 172 1 NR2 $T=366420 920760 0 0 $X=366420 $Y=920380
X4529 160 2 2299 146 1 NR2 $T=368280 920760 0 0 $X=368280 $Y=920380
X4530 169 2 2276 188 1 NR2 $T=370140 930840 0 0 $X=370140 $Y=930460
X4531 186 2 2169 172 1 NR2 $T=371380 900600 0 0 $X=371380 $Y=900220
X4532 187 2 2341 190 1 NR2 $T=373860 900600 0 0 $X=373860 $Y=900220
X4533 97 2 2326 171 1 NR2 $T=373860 910680 1 0 $X=373860 $Y=905260
X4534 160 2 2350 190 1 NR2 $T=373860 920760 0 0 $X=373860 $Y=920380
X4535 113 2 2262 182 1 NR2 $T=373860 940920 0 0 $X=373860 $Y=940540
X4536 118 2 2315 190 1 NR2 $T=377580 910680 0 180 $X=375720 $Y=905260
X4537 2052 2 2327 190 1 NR2 $T=377580 920760 0 180 $X=375720 $Y=915340
X4538 1887 2 2322 171 1 NR2 $T=377580 930840 0 180 $X=375720 $Y=925420
X4539 118 2 2357 146 1 NR2 $T=377580 910680 1 0 $X=377580 $Y=905260
X4540 2052 2 2375 146 1 NR2 $T=380680 920760 0 180 $X=378820 $Y=915340
X4541 2052 2 2366 66 1 NR2 $T=381300 910680 0 180 $X=379440 $Y=905260
X4542 2248 2 2372 200 1 NR2 $T=382540 920760 1 0 $X=382540 $Y=915340
X4543 202 2 199 203 1 NR2 $T=385640 900600 0 0 $X=385640 $Y=900220
X4544 81 2 2363 188 1 NR2 $T=386260 920760 1 0 $X=386260 $Y=915340
X4545 169 2 2352 203 1 NR2 $T=388120 930840 1 180 $X=386260 $Y=930460
X4546 169 2 2447 200 1 NR2 $T=391840 920760 1 0 $X=391840 $Y=915340
X4547 97 2 2475 2215 1 NR2 $T=394940 900600 0 0 $X=394940 $Y=900220
X4548 174 2 2473 200 1 NR2 $T=396800 920760 1 0 $X=396800 $Y=915340
X4549 174 2 2463 188 1 NR2 $T=396800 930840 0 0 $X=396800 $Y=930460
X4550 186 2 2485 2215 1 NR2 $T=400520 900600 1 180 $X=398660 $Y=900220
X4551 2877 2 2879 2723 1 NR2 $T=464380 1071960 0 0 $X=464380 $Y=1071580
X4552 2972 2 2968 2701 1 NR2 $T=482360 1071960 0 180 $X=480500 $Y=1066540
X4553 2981 2 2980 2495 1 NR2 $T=483600 1071960 1 180 $X=481740 $Y=1071580
X4554 3024 2 3035 2553 1 NR2 $T=491040 1061880 0 0 $X=491040 $Y=1061500
X4555 3047 2 3055 2789 1 NR2 $T=496000 1061880 1 180 $X=494140 $Y=1061500
X4556 3033 2 3041 2512 1 NR2 $T=496000 1071960 0 180 $X=494140 $Y=1066540
X4557 3063 2 3075 2849 1 NR2 $T=500960 1041720 0 0 $X=500960 $Y=1041340
X4558 3074 2 3089 2931 1 NR2 $T=503440 1021560 1 0 $X=503440 $Y=1016140
X4559 3087 2 3097 2859 1 NR2 $T=504680 1051800 1 0 $X=504680 $Y=1046380
X4560 3085 2 3088 341 1 NR2 $T=505300 971160 1 0 $X=505300 $Y=965740
X4561 3086 2 3093 342 1 NR2 $T=505300 1001400 1 0 $X=505300 $Y=995980
X4562 347 2 3104 342 1 NR2 $T=510260 940920 0 180 $X=508400 $Y=935500
X4563 3096 2 3095 341 1 NR2 $T=510260 951000 1 180 $X=508400 $Y=950620
X4564 350 2 3122 342 1 NR2 $T=512120 1001400 0 180 $X=510260 $Y=995980
X4565 3120 2 3129 2900 1 NR2 $T=512120 1031640 0 180 $X=510260 $Y=1026220
X4566 3305 2 3301 341 1 NR2 $T=544360 971160 0 180 $X=542500 $Y=965740
X4567 3328 2 3314 341 1 NR2 $T=548080 951000 0 180 $X=546220 $Y=945580
X4568 3085 2 3531 470 1 NR2 $T=585280 971160 1 0 $X=585280 $Y=965740
X4569 3328 2 3584 489 1 NR2 $T=598920 940920 0 0 $X=598920 $Y=940540
X4570 489 2 3606 3305 1 NR2 $T=604500 951000 0 0 $X=604500 $Y=950620
X4571 3681 2 3675 516 1 NR2 $T=615660 1071960 1 180 $X=613800 $Y=1071580
X4572 3671 2 3688 522 1 NR2 $T=616280 1082040 0 0 $X=616280 $Y=1081660
X4573 3701 2 3690 3392 1 NR2 $T=618760 1061880 1 180 $X=616900 $Y=1061500
X4574 3721 2 3715 3424 1 NR2 $T=621860 1061880 1 180 $X=620000 $Y=1061500
X4575 3725 2 3735 533 1 NR2 $T=622480 1051800 1 0 $X=622480 $Y=1046380
X4576 489 2 3739 3085 1 NR2 $T=624960 951000 0 0 $X=624960 $Y=950620
X4577 3096 2 3801 489 1 NR2 $T=639840 951000 0 180 $X=637980 $Y=945580
X4578 3085 2 3951 596 1 NR2 $T=664020 951000 0 0 $X=664020 $Y=950620
X4579 3916 2 3944 3959 1 NR2 $T=664020 1071960 0 0 $X=664020 $Y=1071580
X4580 3962 2 3896 600 1 NR2 $T=667120 961080 1 0 $X=667120 $Y=955660
X4581 3964 2 3968 3486 1 NR2 $T=667120 1021560 1 0 $X=667120 $Y=1016140
X4582 3994 2 3984 600 1 NR2 $T=673320 961080 1 180 $X=671460 $Y=960700
X4583 608 2 3983 596 1 NR2 $T=672700 951000 1 0 $X=672700 $Y=945580
X4584 4030 2 4021 3894 1 NR2 $T=677660 920760 1 180 $X=675800 $Y=920380
X4585 4015 2 4014 350 1 NR2 $T=675800 1001400 1 0 $X=675800 $Y=995980
X4586 4015 2 3914 3086 1 NR2 $T=675800 1001400 0 0 $X=675800 $Y=1001020
X4587 4015 2 3980 3962 1 NR2 $T=680760 1001400 1 0 $X=680760 $Y=995980
X4588 4081 2 4053 3495 1 NR2 $T=682620 1031640 0 180 $X=680760 $Y=1026220
X4589 4062 2 4079 4072 1 NR2 $T=682620 1082040 1 0 $X=682620 $Y=1076620
X4590 4089 2 4093 3287 1 NR2 $T=688200 1041720 1 180 $X=686340 $Y=1041340
X4591 4167 2 4166 3159 1 NR2 $T=700600 1051800 1 180 $X=698740 $Y=1051420
X4592 4279 2 4272 3323 1 NR2 $T=721680 1041720 0 180 $X=719820 $Y=1036300
X4593 4288 2 4281 600 1 NR2 $T=724160 951000 0 0 $X=724160 $Y=950620
X4594 4324 2 4322 600 1 NR2 $T=728500 951000 1 180 $X=726640 $Y=950620
X4595 4255 2 4329 4316 1 NR2 $T=727260 1082040 1 0 $X=727260 $Y=1076620
X4596 4339 2 4336 3266 1 NR2 $T=730980 1051800 1 180 $X=729120 $Y=1051420
X4597 4269 2 4349 4350 1 NR2 $T=729120 1082040 1 0 $X=729120 $Y=1076620
X4598 4367 2 4361 3158 1 NR2 $T=734080 1051800 0 180 $X=732220 $Y=1046380
X4599 4360 2 4362 3221 1 NR2 $T=734080 1061880 0 180 $X=732220 $Y=1056460
X4600 347 2 4418 4015 1 NR2 $T=744000 991320 0 180 $X=742140 $Y=985900
X4601 4324 2 4601 4611 1 NR2 $T=775620 971160 0 0 $X=775620 $Y=970780
X4602 4324 2 4792 759 1 NR2 $T=804140 981240 0 0 $X=804140 $Y=980860
X4603 4288 2 4852 831 1 NR2 $T=812820 1011480 1 0 $X=812820 $Y=1006060
X4604 4896 2 4890 831 1 NR2 $T=820880 1001400 0 180 $X=819020 $Y=995980
X4605 718 2 4926 3994 1 NR2 $T=826460 951000 1 0 $X=826460 $Y=945580
X4606 347 2 4927 4611 1 NR2 $T=827080 961080 0 0 $X=827080 $Y=960700
X4607 350 2 4990 831 1 NR2 $T=838860 1001400 1 0 $X=838860 $Y=995980
X4608 5009 2 5006 3962 1 NR2 $T=843200 1001400 0 180 $X=841340 $Y=995980
X4609 5009 2 5027 3086 1 NR2 $T=844440 981240 1 0 $X=844440 $Y=975820
X4610 3962 2 5029 831 1 NR2 $T=846300 1001400 0 180 $X=844440 $Y=995980
X4611 5009 2 5041 3994 1 NR2 $T=846300 1001400 1 0 $X=846300 $Y=995980
X4612 872 2 5098 5020 1 NR2 $T=855600 940920 0 0 $X=855600 $Y=940540
X4613 3994 2 5249 759 1 NR2 $T=882880 991320 1 180 $X=881020 $Y=990940
X4614 3962 2 5270 759 1 NR2 $T=883500 1001400 1 180 $X=881640 $Y=1001020
X4615 5460 2 3976 978 1 NR2 $T=921940 951000 1 180 $X=920080 $Y=950620
X4616 347 2 5454 5463 1 NR2 $T=920700 951000 1 0 $X=920700 $Y=945580
X4617 4324 2 5485 5463 1 NR2 $T=923180 951000 1 0 $X=923180 $Y=945580
X4618 3994 2 5499 5463 1 NR2 $T=925660 951000 0 0 $X=925660 $Y=950620
X4619 3086 2 5533 5463 1 NR2 $T=928760 951000 0 0 $X=928760 $Y=950620
X4620 4896 2 5535 5463 1 NR2 $T=933720 940920 0 0 $X=933720 $Y=940540
X4621 5577 2 5572 993 1 NR2 $T=940540 940920 0 180 $X=938680 $Y=935500
X4622 5020 2 5663 5463 1 NR2 $T=952940 940920 0 180 $X=951080 $Y=935500
X4623 4896 2 5907 1097 1 NR2 $T=1001920 940920 1 0 $X=1001920 $Y=935500
X4624 4896 2 6050 1150 1 NR2 $T=1029200 951000 1 0 $X=1029200 $Y=945580
X4625 4896 2 6075 1157 1 NR2 $T=1031060 951000 1 0 $X=1031060 $Y=945580
X4626 5577 2 6188 1097 1 NR2 $T=1054000 940920 0 180 $X=1052140 $Y=935500
X4627 5577 2 6185 1150 1 NR2 $T=1054000 951000 1 0 $X=1054000 $Y=945580
X4628 5020 2 6196 1150 1 NR2 $T=1057720 951000 0 180 $X=1055860 $Y=945580
X4629 5020 2 6211 1157 1 NR2 $T=1057720 951000 1 0 $X=1057720 $Y=945580
X4630 5577 2 6200 1157 1 NR2 $T=1057720 951000 0 0 $X=1057720 $Y=950620
X4631 2298 4 1 2 INV12CK $T=369520 1051800 0 180 $X=359600 $Y=1046380
X4632 2298 185 1 2 INV12CK $T=383160 1051800 0 180 $X=373240 $Y=1046380
X4633 318 2637 1 2 INV12CK $T=489180 940920 0 180 $X=479260 $Y=935500
X4634 318 253 1 2 INV12CK $T=490420 920760 0 180 $X=480500 $Y=915340
X4635 3056 252 1 2 INV12CK $T=506540 1031640 0 180 $X=496620 $Y=1026220
X4636 3056 3257 1 2 INV12CK $T=546220 1041720 0 180 $X=536300 $Y=1036300
X4637 3056 399 1 2 INV12CK $T=546840 1051800 0 0 $X=546840 $Y=1051420
X4638 247 3673 1 2 INV12CK $T=607600 961080 0 0 $X=607600 $Y=960700
X4639 3768 380 1 2 INV12CK $T=629300 971160 0 0 $X=629300 $Y=970780
X4640 576 3768 1 2 INV12CK $T=652860 971160 0 0 $X=652860 $Y=970780
X4641 3768 3819 1 2 INV12CK $T=698120 971160 0 180 $X=688200 $Y=965740
X4642 3768 4341 1 2 INV12CK $T=755780 971160 0 0 $X=755780 $Y=970780
X4643 4687 599 1 2 INV12CK $T=789880 1041720 0 180 $X=779960 $Y=1036300
X4644 4687 799 1 2 INV12CK $T=809100 1031640 0 0 $X=809100 $Y=1031260
X4645 4687 4870 1 2 INV12CK $T=811580 1021560 0 0 $X=811580 $Y=1021180
X4646 5711 946 1 2 INV12CK $T=966580 1051800 0 180 $X=956660 $Y=1046380
X4647 5711 5328 1 2 INV12CK $T=962240 1011480 1 0 $X=962240 $Y=1006060
X4648 5964 6041 1 2 INV12CK $T=1067020 1011480 0 0 $X=1067020 $Y=1011100
X4649 5964 1149 1 2 INV12CK $T=1076320 1071960 0 0 $X=1076320 $Y=1071580
X4650 141 130 2 1 2019 OR2 $T=338520 1082040 1 180 $X=336040 $Y=1081660
X4651 336 3085 2 1 2838 OR2 $T=505300 981240 0 180 $X=502820 $Y=975820
X4652 336 3086 2 1 2947 OR2 $T=505300 981240 1 180 $X=502820 $Y=980860
X4653 336 3096 2 1 2945 OR2 $T=507160 961080 1 180 $X=504680 $Y=960700
X4654 342 346 2 1 2744 OR2 $T=509020 961080 0 180 $X=506540 $Y=955660
X4655 336 347 2 1 2948 OR2 $T=510880 961080 1 180 $X=508400 $Y=960700
X4656 373 3085 2 1 3169 OR2 $T=531960 971160 0 180 $X=529480 $Y=965740
X4657 373 3096 2 1 3222 OR2 $T=536920 951000 1 0 $X=536920 $Y=945580
X4658 373 3305 2 1 3321 OR2 $T=544980 971160 0 0 $X=544980 $Y=970780
X4659 373 3328 2 1 3343 OR2 $T=553660 951000 0 180 $X=551180 $Y=945580
X4660 470 3096 2 1 3440 OR2 $T=584660 961080 1 180 $X=582180 $Y=960700
X4661 470 3328 2 1 3414 OR2 $T=585280 940920 0 0 $X=585280 $Y=940540
X4662 470 3305 2 1 3558 OR2 $T=599540 971160 0 180 $X=597060 $Y=965740
X4663 596 3096 2 1 4164 OR2 $T=702460 951000 0 180 $X=699980 $Y=945580
X4664 596 4263 2 1 4227 OR2 $T=717960 940920 0 0 $X=717960 $Y=940540
X4665 4015 4288 2 1 4353 OR2 $T=730360 991320 0 0 $X=730360 $Y=990940
X4666 4015 346 2 1 4381 OR2 $T=745240 961080 1 180 $X=742760 $Y=960700
X4667 718 4324 2 1 4446 OR2 $T=748340 961080 0 0 $X=748340 $Y=960700
X4668 759 4288 2 1 4532 OR2 $T=775620 1001400 1 180 $X=773140 $Y=1001020
X4669 4611 346 2 1 4539 OR2 $T=777480 961080 1 180 $X=775000 $Y=960700
X4670 4611 4288 2 1 4695 OR2 $T=805380 971160 1 180 $X=802900 $Y=970780
X4671 5402 5474 2 1 5460 OR2 $T=924420 951000 1 180 $X=921940 $Y=950620
X4672 1080 4896 2 1 5828 OR2 $T=990760 940920 0 180 $X=988280 $Y=935500
X4673 1080 4263 2 1 5856 OR2 $T=995100 940920 1 0 $X=995100 $Y=935500
X4674 1097 4263 2 1 5930 OR2 $T=1005640 940920 1 0 $X=1005640 $Y=935500
X4675 1150 4263 2 1 6000 OR2 $T=1026100 940920 1 180 $X=1023620 $Y=940540
X4676 1080 5020 2 1 6088 OR2 $T=1037260 940920 1 0 $X=1037260 $Y=935500
X4677 1157 4263 2 1 6119 OR2 $T=1037880 951000 1 0 $X=1037880 $Y=945580
X4678 1080 5577 2 1 6125 OR2 $T=1039740 940920 1 0 $X=1039740 $Y=935500
X4679 1097 5020 2 1 6186 OR2 $T=1052140 930840 0 0 $X=1052140 $Y=930460
X4680 1632 1619 1595 1636 2 1 1557 OA22 $T=274040 930840 0 180 $X=269700 $Y=925420
X4681 1762 1777 1742 1763 2 1 1781 OA22 $T=289540 940920 1 0 $X=289540 $Y=935500
X4682 1652 1776 1785 1769 2 1 1773 OA22 $T=294500 1041720 0 180 $X=290160 $Y=1036300
X4683 192 2209 2323 2358 2 1 2386 OA22 $T=379440 951000 1 0 $X=379440 $Y=945580
X4684 14 1403 1 2 1393 AN2 $T=234360 1031640 0 0 $X=234360 $Y=1031260
X4685 1333 1386 1 2 1430 AN2 $T=241800 1031640 0 180 $X=239320 $Y=1026220
X4686 1452 1417 1 2 1441 AN2 $T=242420 1051800 0 180 $X=239940 $Y=1046380
X4687 34 1541 1 2 1506 AN2 $T=256680 1021560 0 180 $X=254200 $Y=1016140
X4688 1516 1558 1 2 1552 AN2 $T=257920 961080 1 0 $X=257920 $Y=955660
X4689 40 1609 1 2 1448 AN2 $T=266600 1031640 1 180 $X=264120 $Y=1031260
X4690 1640 1448 1 2 1613 AN2 $T=270320 1041720 0 180 $X=267840 $Y=1036300
X4691 1659 1656 1 2 1628 AN2 $T=272800 961080 1 180 $X=270320 $Y=960700
X4692 1538 1609 1 2 1792 AN2 $T=289540 1041720 0 0 $X=289540 $Y=1041340
X4693 1947 1961 1 2 1967 AN2 $T=316820 971160 1 0 $X=316820 $Y=965740
X4694 1960 1993 1 2 2004 AN2 $T=323640 961080 1 0 $X=323640 $Y=955660
X4695 2045 2048 1 2 2072 AN2 $T=332320 971160 1 0 $X=332320 $Y=965740
X4696 2027 2079 1 2 2054 AN2 $T=336660 1071960 1 180 $X=334180 $Y=1071580
X4697 2015 2092 1 2 2125 AN2 $T=340380 961080 1 0 $X=340380 $Y=955660
X4698 4644 4631 1 2 768 AN2 $T=782440 1051800 0 180 $X=779960 $Y=1046380
X4699 1953 2 2019 1957 91 1 NR3 $T=323640 1082040 1 0 $X=323640 $Y=1076620
X4700 2098 2 2109 2115 147 1 NR3 $T=338520 1061880 0 0 $X=338520 $Y=1061500
X4701 783 2 4685 4690 4657 1 NR3 $T=788020 1061880 1 0 $X=788020 $Y=1056460
X4702 4706 2 4702 4705 4638 1 NR3 $T=791120 1011480 0 0 $X=791120 $Y=1011100
X4703 794 2 4675 4723 4672 1 NR3 $T=792360 1061880 1 0 $X=792360 $Y=1056460
X4704 800 2 4720 4732 4694 1 NR3 $T=794220 1041720 1 0 $X=794220 $Y=1036300
X4705 4741 2 4736 4758 4716 1 NR3 $T=797320 1051800 0 0 $X=797320 $Y=1051420
X4706 4743 2 4738 814 4735 1 NR3 $T=798560 1071960 1 0 $X=798560 $Y=1066540
X4707 816 2 4788 4790 4652 1 NR3 $T=802900 1041720 1 0 $X=802900 $Y=1036300
X4708 837 2 4869 4868 4050 1 NR3 $T=817160 961080 1 180 $X=814060 $Y=960700
X4709 840 2 4878 4825 4304 1 NR3 $T=818400 930840 1 180 $X=815300 $Y=930460
X4710 845 2 4885 4838 4047 1 NR3 $T=820260 940920 1 180 $X=817160 $Y=940540
X4711 849 2 4907 4905 4264 1 NR3 $T=823980 971160 0 180 $X=820880 $Y=965740
X4712 873 2 5026 4893 4190 1 NR3 $T=846300 951000 1 180 $X=843200 $Y=950620
X4713 875 2 4998 5052 4858 1 NR3 $T=846920 1071960 1 0 $X=846920 $Y=1066540
X4714 878 2 4984 5058 4826 1 NR3 $T=848160 1031640 1 0 $X=848160 $Y=1026220
X4715 5125 2 5057 5131 4749 1 NR3 $T=861180 1061880 0 0 $X=861180 $Y=1061500
X4716 904 2 5144 5169 4752 1 NR3 $T=866760 1051800 1 0 $X=866760 $Y=1046380
X4717 5168 2 5166 5174 4843 1 NR3 $T=867380 1031640 0 0 $X=867380 $Y=1031260
X4718 5198 2 5206 5212 4765 1 NR3 $T=873580 1001400 0 0 $X=873580 $Y=1001020
X4719 955 2 5374 5357 3996 1 NR3 $T=903340 971160 0 180 $X=900240 $Y=965740
X4720 985 2 5461 5403 3946 1 NR3 $T=923800 971160 1 180 $X=920700 $Y=970780
X4721 983 2 5475 5369 3995 1 NR3 $T=921940 961080 1 0 $X=921940 $Y=955660
X4722 1449 1439 1 1423 2 OR2B1S $T=243660 1082040 1 0 $X=243660 $Y=1076620
X4723 2174 2198 1 2244 2 OR2B1S $T=358980 1031640 1 0 $X=358980 $Y=1026220
X4724 2805 2799 1 2759 2 OR2B1S $T=452600 1001400 1 180 $X=449500 $Y=1001020
X4725 2906 2925 1 2940 2 OR2B1S $T=474920 940920 0 0 $X=474920 $Y=940540
X4726 5223 5435 1 5429 2 OR2B1S $T=919460 940920 1 180 $X=916360 $Y=940540
X4727 2470 2385 2 1 2494 218 2446 208 2455 2292 2440 1299 ICV_7 $T=392460 1071960 1 0 $X=392460 $Y=1066540
X4728 2822 2385 2 1 2893 2819 2728 2483 2855 2740 2798 1299 ICV_7 $T=460040 1061880 1 0 $X=460040 $Y=1056460
X4729 3000 2993 2 1 2923 3023 2710 2979 2937 2986 2987 1299 ICV_7 $T=482980 1001400 0 0 $X=482980 $Y=1001020
X4730 2575 2945 2 1 2946 3062 2579 2884 3025 2222 2548 1299 ICV_7 $T=491040 971160 1 0 $X=491040 $Y=965740
X4731 3536 3417 2 1 3554 3548 3396 3400 465 467 3527 1299 ICV_7 $T=582180 1082040 1 0 $X=582180 $Y=1076620
X4732 3769 3682 2 1 3793 3747 3674 3656 3731 3744 3743 1299 ICV_7 $T=624960 1051800 0 0 $X=624960 $Y=1051420
X4733 3931 3682 2 1 3967 3969 3836 3832 3911 3919 3923 1299 ICV_7 $T=657820 1051800 1 0 $X=657820 $Y=1046380
X4734 3925 4080 2 1 4101 607 3999 3961 4059 3851 3954 1299 ICV_7 $T=681380 940920 0 0 $X=681380 $Y=940540
X4735 4094 634 2 1 4109 3722 626 601 4074 624 4076 1299 ICV_7 $T=683860 910680 1 0 $X=683860 $Y=905260
X4736 4398 4061 2 1 4410 709 4315 4100 4363 4386 4337 1299 ICV_7 $T=735320 1061880 0 0 $X=735320 $Y=1061500
X4737 764 4505 2 1 4643 4635 4576 4540 4590 4463 762 1299 ICV_7 $T=774380 971160 1 0 $X=774380 $Y=965740
X4738 5797 5796 2 1 5822 5594 5707 5548 5780 1068 5785 1299 ICV_7 $T=976500 940920 1 0 $X=976500 $Y=935500
X4739 6059 1151 2 1 6068 5809 1148 1140 5971 6055 6022 1299 ICV_7 $T=1024860 1061880 0 0 $X=1024860 $Y=1061500
X4740 6133 1169 2 1 6163 5976 6108 6113 5940 5980 6124 1299 ICV_7 $T=1038500 1041720 1 0 $X=1038500 $Y=1036300
X4741 6478 6415 2 1 6495 6366 6440 1247 6431 6461 6439 1299 ICV_7 $T=1107320 951000 1 0 $X=1107320 $Y=945580
X4742 6502 6408 2 1 6521 6366 6223 1173 6435 6505 6509 1299 ICV_7 $T=1116000 951000 0 0 $X=1116000 $Y=950620
X4743 2658 1 2 2683 2741 252 2614 248 1299 ICV_8 $T=425320 1041720 0 0 $X=425320 $Y=1041340
X4744 3029 1 2 3052 3090 252 309 3029 1299 ICV_8 $T=491660 1082040 0 0 $X=491660 $Y=1081660
X4745 3269 1 2 3292 3338 3257 3306 3269 1299 ICV_8 $T=537540 1041720 0 0 $X=537540 $Y=1041340
X4746 3324 1 2 3351 3403 3257 3307 3324 1299 ICV_8 $T=547460 991320 1 0 $X=547460 $Y=985900
X4747 3825 1 2 3845 3885 3819 3821 3643 1299 ICV_8 $T=642940 930840 0 0 $X=642940 $Y=930460
X4748 3907 1 2 3933 3998 3819 3901 3563 1299 ICV_8 $T=658440 991320 1 0 $X=658440 $Y=985900
X4749 3918 1 2 3943 4004 3819 3972 3918 1299 ICV_8 $T=659680 1021560 0 0 $X=659680 $Y=1021180
X4750 4784 1 2 4819 4836 4870 4778 4733 1299 ICV_8 $T=803520 991320 0 0 $X=803520 $Y=990940
X4751 4972 1 2 4999 5075 4870 4935 5015 1299 ICV_8 $T=838240 971160 0 0 $X=838240 $Y=970780
X4752 5521 1 2 5513 5568 973 5589 5573 1299 ICV_8 $T=934960 951000 1 0 $X=934960 $Y=945580
X4753 5756 1 2 5775 5802 5328 5697 5756 1299 ICV_8 $T=970920 991320 1 0 $X=970920 $Y=985900
X4754 5841 1 2 5894 6001 946 1118 5941 1299 ICV_8 $T=1001920 1061880 1 0 $X=1001920 $Y=1056460
X4755 5941 1 2 5998 5993 946 1135 1111 1299 ICV_8 $T=1014320 1071960 0 0 $X=1014320 $Y=1071580
X4756 5980 1 2 6016 6034 1149 5910 6015 1299 ICV_8 $T=1014940 1051800 1 0 $X=1014940 $Y=1046380
X4757 5996 1 2 6072 6184 6041 6126 6122 1299 ICV_8 $T=1039740 981240 0 0 $X=1039740 $Y=980860
X4758 6118 1 2 6127 6151 1149 6093 6118 1299 ICV_8 $T=1039740 1031640 1 0 $X=1039740 $Y=1026220
X4759 6220 1 2 6253 6297 1149 6236 6257 1299 ICV_8 $T=1061440 1061880 0 0 $X=1061440 $Y=1061500
X4760 6143 1 2 6155 6217 6041 6162 6232 1299 ICV_8 $T=1065160 961080 0 0 $X=1065160 $Y=960700
X4761 6291 1 2 6309 6365 1149 6194 6311 1299 ICV_8 $T=1075080 1031640 1 0 $X=1075080 $Y=1026220
X4762 6482 1 2 6491 6517 1149 6450 6447 1299 ICV_8 $T=1112280 1031640 1 0 $X=1112280 $Y=1026220
X4763 6460 1 2 6484 6499 1149 6512 6446 1299 ICV_8 $T=1112280 1061880 1 0 $X=1112280 $Y=1056460
X4764 303 2385 2 1 2952 2888 2908 2904 2854 300 301 1299 ICV_9 $T=470580 1031640 0 0 $X=470580 $Y=1031260
X4765 3296 3195 2 1 3320 339 3185 3192 3270 3260 381 1299 ICV_9 $T=538780 1061880 0 0 $X=538780 $Y=1061500
X4766 3382 3378 2 1 3404 3217 3311 3293 3282 3324 3355 1299 ICV_9 $T=553660 981240 0 0 $X=553660 $Y=980860
X4767 2653 482 2 1 3613 3556 484 413 3564 487 3589 1299 ICV_9 $T=597060 920760 0 0 $X=597060 $Y=920380
X4768 3912 3682 2 1 3936 3863 3836 3832 3897 3899 3908 1299 ICV_9 $T=655340 1061880 1 0 $X=655340 $Y=1056460
X4769 4318 4149 2 1 4344 3806 4278 4271 4290 4195 4277 1299 ICV_9 $T=722920 1031640 1 0 $X=722920 $Y=1026220
X4770 4295 3975 2 1 4352 485 3999 3961 4302 687 4270 1299 ICV_9 $T=724160 940920 0 0 $X=724160 $Y=940540
X4771 4369 4149 2 1 4407 4378 4278 4271 4346 4356 697 1299 ICV_9 $T=730360 1031640 0 0 $X=730360 $Y=1031260
X4772 4389 4061 2 1 4406 4378 4315 4100 4355 4377 4376 1299 ICV_9 $T=733460 1051800 0 0 $X=733460 $Y=1051420
X4773 4919 4923 2 1 4938 4131 4848 823 4747 848 4915 1299 ICV_9 $T=821500 1071960 1 0 $X=821500 $Y=1066540
X4774 900 4933 2 1 5164 5070 4959 4995 5120 4960 896 1299 ICV_9 $T=860560 920760 1 0 $X=860560 $Y=915340
X4775 5291 917 2 1 5319 868 923 925 5181 5276 928 1299 ICV_9 $T=883500 1082040 0 0 $X=883500 $Y=1081660
X4776 996 5452 2 1 5411 971 5465 5453 5482 5424 994 1299 ICV_9 $T=923800 1061880 0 0 $X=923800 $Y=1061500
X4777 5543 5452 2 1 5564 5575 5465 5453 1006 1008 5501 1299 ICV_9 $T=931860 1061880 0 0 $X=931860 $Y=1061500
X4778 5605 5609 2 1 5634 5618 1021 5548 5585 5491 5590 1299 ICV_9 $T=941780 930840 0 0 $X=941780 $Y=930460
X4779 5692 5678 2 1 5715 5598 5654 5646 5670 5658 5684 1299 ICV_9 $T=955420 1011480 0 0 $X=955420 $Y=1011100
X4780 1058 5657 2 1 5753 5433 5655 5644 5701 1053 5725 1299 ICV_9 $T=962860 1061880 0 0 $X=962860 $Y=1061500
X4781 5739 5627 2 1 5755 971 5655 5644 5712 5734 5702 1299 ICV_9 $T=964100 1041720 1 0 $X=964100 $Y=1036300
X4782 5784 5779 2 1 5794 5729 5553 1052 5751 5767 5768 1299 ICV_9 $T=972780 981240 1 0 $X=972780 $Y=975820
X4783 5999 5986 2 1 5927 6024 5962 5937 5969 5985 1131 1299 ICV_9 $T=1013700 1001400 1 0 $X=1013700 $Y=995980
X4784 6127 6116 2 1 6151 5900 6108 6113 5923 6118 1164 1299 ICV_9 $T=1037880 1021560 0 0 $X=1037880 $Y=1021180
X4785 6152 1160 2 1 6172 1176 1168 1165 5942 6128 6073 1299 ICV_9 $T=1042840 1071960 0 0 $X=1042840 $Y=1071580
X4786 6470 1268 2 1 6494 1238 1256 6412 6454 6460 6463 1299 ICV_9 $T=1106700 1082040 1 0 $X=1106700 $Y=1076620
X4787 6474 1193 2 1 6489 1279 1260 6348 1270 6433 1275 1299 ICV_9 $T=1107320 900600 0 0 $X=1107320 $Y=900220
X4788 6480 1268 2 1 6508 6330 6416 6304 6407 6471 6447 1299 ICV_9 $T=1108560 1021560 1 0 $X=1108560 $Y=1016140
X4789 6491 6486 2 1 6511 6442 6416 6304 6403 6487 6482 1299 ICV_9 $T=1109800 1031640 0 0 $X=1109800 $Y=1031260
X4790 2620 1 2 2649 2685 185 2614 2620 1299 ICV_10 $T=431520 1061880 0 180 $X=419740 $Y=1056460
X4791 2704 1 2 2688 2633 2637 2651 2477 1299 ICV_10 $T=434000 981240 0 180 $X=422220 $Y=975820
X4792 2667 1 2 2751 2733 2637 2644 2676 1299 ICV_10 $T=440200 1021560 0 180 $X=428420 $Y=1016140
X4793 2757 1 2 2777 2845 2637 2734 2795 1299 ICV_10 $T=461280 1001400 0 180 $X=449500 $Y=995980
X4794 2853 1 2 2836 2858 253 2753 2532 1299 ICV_10 $T=463140 930840 1 180 $X=451360 $Y=930460
X4795 2862 1 2 2878 2895 253 279 2862 1299 ICV_10 $T=474300 910680 1 180 $X=462520 $Y=910300
X4796 2987 1 2 3000 3061 2637 2887 2985 1299 ICV_10 $T=500340 1011480 0 180 $X=488560 $Y=1006060
X4797 3171 1 2 3201 3135 252 3079 3100 1299 ICV_10 $T=519560 1041720 0 180 $X=507780 $Y=1036300
X4798 3544 1 2 3565 3525 3257 3473 437 1299 ICV_10 $T=591480 981240 0 180 $X=579700 $Y=975820
X4799 3521 1 2 3513 3580 380 3461 3520 1299 ICV_10 $T=600160 910680 1 180 $X=588380 $Y=910300
X4800 3869 1 2 3866 3857 3819 3794 553 1299 ICV_10 $T=651620 981240 1 180 $X=639840 $Y=980860
X4801 4364 1 2 4397 4390 599 4268 4321 1299 ICV_10 $T=739040 1071960 1 180 $X=727260 $Y=1071580
X4802 4448 1 2 4477 4422 4341 4332 3577 1299 ICV_10 $T=750820 971160 1 180 $X=739040 $Y=970780
X4803 693 1 2 737 4494 686 717 719 1299 ICV_10 $T=761360 900600 1 180 $X=749580 $Y=900220
X4804 4937 1 2 4973 4991 4870 4942 4937 1299 ICV_10 $T=840720 1021560 0 180 $X=828940 $Y=1016140
X4805 892 1 2 5089 5097 799 862 874 1299 ICV_10 $T=857460 1082040 0 180 $X=845680 $Y=1076620
X4806 5047 1 2 5102 5106 799 5064 5047 1299 ICV_10 $T=859320 1061880 0 180 $X=847540 $Y=1056460
X4807 5370 1 2 5388 5394 869 5399 949 1299 ICV_10 $T=915740 930840 1 180 $X=903960 $Y=930460
X4808 5569 1 2 5613 5748 973 5682 5691 1299 ICV_10 $T=970920 940920 1 180 $X=959140 $Y=940540
X4809 5734 1 2 5761 5755 5328 5717 5702 1299 ICV_10 $T=972160 1031640 0 180 $X=960380 $Y=1026220
X4810 5786 1 2 5750 1073 973 1023 5736 1299 ICV_10 $T=982080 900600 1 180 $X=970300 $Y=900220
X4811 5660 1 2 5665 5822 973 5790 5785 1299 ICV_10 $T=988900 930840 0 180 $X=977120 $Y=925420
X4812 5791 1 2 5840 5849 5328 5804 5805 1299 ICV_10 $T=993860 1021560 1 180 $X=982080 $Y=1021180
X4813 6132 1 2 6123 6106 6041 6020 6035 1299 ICV_10 $T=1042840 1011480 0 180 $X=1031060 $Y=1006060
X4814 6055 1 2 6102 6120 1149 5910 6055 1299 ICV_10 $T=1045940 1061880 0 180 $X=1034160 $Y=1056460
X4815 6328 1 2 6384 6456 6041 6346 6411 1299 ICV_10 $T=1109800 1011480 1 180 $X=1098020 $Y=1011100
X4816 2300 1 2 2333 2340 185 2379 2406 1299 ICV_11 $T=370140 1041720 1 0 $X=370140 $Y=1036300
X4817 2305 1 2 2339 2346 185 2380 2256 1299 ICV_11 $T=370760 1011480 1 0 $X=370760 $Y=1006060
X4818 2502 1 2 2536 2546 185 236 2571 1299 ICV_11 $T=403000 1082040 1 0 $X=403000 $Y=1076620
X4819 2516 1 2 2585 2603 185 2651 2639 1299 ICV_11 $T=411680 991320 1 0 $X=411680 $Y=985900
X4820 2795 1 2 2827 2847 2637 2887 2880 1299 ICV_11 $T=453840 1011480 1 0 $X=453840 $Y=1006060
X4821 2872 1 2 2918 2934 252 2950 2996 1299 ICV_11 $T=469960 1041720 1 0 $X=469960 $Y=1036300
X4822 3100 1 2 3116 3161 252 3071 3235 1299 ICV_11 $T=512740 1041720 0 0 $X=512740 $Y=1041340
X4823 3160 1 2 3187 3193 252 372 3250 1299 ICV_11 $T=517700 1082040 1 0 $X=517700 $Y=1076620
X4824 371 1 2 385 3262 252 396 382 1299 ICV_11 $T=531340 1082040 0 0 $X=531340 $Y=1081660
X4825 3499 1 2 3506 3537 3257 3559 3524 1299 ICV_11 $T=580940 1031640 0 0 $X=580940 $Y=1031260
X4826 3507 1 2 3540 3553 399 3592 3570 1299 ICV_11 $T=586520 1061880 1 0 $X=586520 $Y=1056460
X4827 3724 1 2 3734 3760 380 3794 552 1299 ICV_11 $T=621860 971160 1 0 $X=621860 $Y=965740
X4828 4051 1 2 4104 4196 3819 4236 4195 1299 ICV_11 $T=699360 1031640 1 0 $X=699360 $Y=1026220
X4829 4225 1 2 4209 4276 599 4124 4323 1299 ICV_11 $T=715480 1051800 1 0 $X=715480 $Y=1046380
X4830 4425 1 2 4450 4449 4341 4459 4425 1299 ICV_11 $T=745860 1001400 0 0 $X=745860 $Y=1001020
X4831 4460 1 2 4496 4495 4341 4476 4560 1299 ICV_11 $T=754540 920760 0 0 $X=754540 $Y=920380
X4832 4628 1 2 4658 4666 4341 4719 4628 1299 ICV_11 $T=781200 920760 0 0 $X=781200 $Y=920380
X4833 4632 1 2 4665 4671 4341 4692 4632 1299 ICV_11 $T=781820 961080 1 0 $X=781820 $Y=955660
X4834 4751 1 2 4779 4770 4341 4708 4751 1299 ICV_11 $T=797940 1011480 0 0 $X=797940 $Y=1011100
X4835 5710 1 2 5726 5740 973 5682 1067 1299 ICV_11 $T=962240 930840 0 0 $X=962240 $Y=930460
X4836 5785 1 2 5797 5817 973 5790 1088 1299 ICV_11 $T=980220 930840 0 0 $X=980220 $Y=930460
X4837 5924 1 2 5933 5955 946 1135 5934 1299 ICV_11 $T=1005020 1071960 1 0 $X=1005020 $Y=1066540
X4838 1201 1 2 1208 6254 1115 1212 6246 1299 ICV_11 $T=1060820 920760 1 0 $X=1060820 $Y=915340
X4839 1215 1 2 6317 6324 1149 1235 6339 1299 ICV_11 $T=1076320 1082040 0 0 $X=1076320 $Y=1081660
X4840 6371 1 2 6393 6404 6041 6398 1255 1299 ICV_11 $T=1091820 991320 1 0 $X=1091820 $Y=985900
X4841 184 2 2258 1 2294 185 2258 197 1299 ICV_12 $T=367660 1082040 0 0 $X=367660 $Y=1081660
X4842 2332 2 191 1 2296 185 2394 2332 1299 ICV_12 $T=375100 1001400 1 0 $X=375100 $Y=995980
X4843 2373 2 2379 1 2387 185 2379 2349 1299 ICV_12 $T=381300 1031640 0 0 $X=381300 $Y=1031260
X4844 2488 2 231 1 2552 185 2614 2528 1299 ICV_12 $T=409820 1061880 0 0 $X=409820 $Y=1061500
X4845 2838 2 2750 1 2844 2637 2825 2830 1299 ICV_12 $T=457560 981240 0 0 $X=457560 $Y=980860
X4846 4627 2 4482 1 4646 599 4482 4724 1299 ICV_12 $T=781820 1061880 0 0 $X=781820 $Y=1061500
X4847 4696 2 4815 1 4835 799 4766 844 1299 ICV_12 $T=807860 1041720 1 0 $X=807860 $Y=1036300
X4848 775 2 4854 1 4851 686 4908 846 1299 ICV_12 $T=812820 940920 1 0 $X=812820 $Y=935500
X4849 5029 2 5032 1 5040 4870 5063 5051 1299 ICV_12 $T=845060 1001400 0 0 $X=845060 $Y=1001020
X4850 5046 2 5055 1 5090 799 5132 902 1299 ICV_12 $T=853740 1031640 1 0 $X=853740 $Y=1026220
X4851 5270 2 5269 1 5283 4870 5333 5259 1299 ICV_12 $T=884740 1001400 0 0 $X=884740 $Y=1001020
X4852 5454 2 5457 1 5468 973 5446 5521 1299 ICV_12 $T=920700 940920 0 0 $X=920700 $Y=940540
X4853 5764 2 5809 1 5816 946 1076 5868 1299 ICV_12 $T=983320 1071960 1 0 $X=983320 $Y=1066540
X4854 5182 2 5847 1 5881 5328 5847 5884 1299 ICV_12 $T=996960 1031640 0 0 $X=996960 $Y=1031260
X4855 1137 2 6076 1 6084 6041 6029 1171 1299 ICV_12 $T=1032300 961080 1 0 $X=1032300 $Y=955660
X4856 6188 2 6197 1 6198 6041 6146 6244 1299 ICV_12 $T=1055860 940920 1 0 $X=1055860 $Y=935500
X4857 1161 2 6261 1 6268 1115 1214 6159 1299 ICV_12 $T=1067020 910680 0 0 $X=1067020 $Y=910300
X4858 6354 2 6363 1 6367 6041 6363 6381 1299 ICV_12 $T=1089340 951000 0 0 $X=1089340 $Y=950620
X4859 204 205 2 1 2294 198 211 208 2434 207 197 1299 ICV_13 $T=386880 1082040 1 180 $X=382540 $Y=1081660
X4860 2415 2398 2 1 2277 193 2433 2419 209 2390 2356 1299 ICV_13 $T=387500 1051800 0 180 $X=383160 $Y=1046380
X4861 2416 2420 2 1 2303 193 2446 208 2428 2381 2355 1299 ICV_13 $T=388120 1071960 0 180 $X=383780 $Y=1066540
X4862 2510 2517 2 1 2441 2488 2539 2523 2531 2516 2383 1299 ICV_13 $T=403620 1001400 1 180 $X=399280 $Y=1001020
X4863 2663 2411 2 1 2630 241 2680 2556 2673 2668 2667 1299 ICV_13 $T=425940 1051800 0 180 $X=421600 $Y=1046380
X4864 2751 2549 2 1 2707 241 2680 2556 2779 2709 248 1299 ICV_13 $T=443920 1051800 0 180 $X=439580 $Y=1046380
X4865 283 260 2 1 278 277 289 286 291 281 2717 1299 ICV_13 $T=458800 900600 1 180 $X=454460 $Y=900220
X4866 3347 3343 2 1 3281 3067 3364 413 3319 3339 409 1299 ICV_13 $T=551180 951000 1 180 $X=546840 $Y=950620
X4867 3361 412 2 1 404 402 387 384 3387 410 416 1299 ICV_13 $T=553660 1082040 1 180 $X=549320 $Y=1081660
X4868 3367 3358 2 1 3335 2902 415 403 3381 3275 3370 1299 ICV_13 $T=554900 920760 1 180 $X=550560 $Y=920380
X4869 3513 455 2 1 3493 294 473 469 3498 3521 3520 1299 ICV_13 $T=583420 910680 1 180 $X=579080 $Y=910300
X4870 3600 3644 2 1 3557 501 3674 3656 3678 3570 3612 1299 ICV_13 $T=613180 1051800 1 180 $X=608840 $Y=1051420
X4871 3729 3746 2 1 3703 3654 3758 3748 3751 3650 3638 1299 ICV_13 $T=623720 991320 0 180 $X=619380 $Y=985900
X4872 3822 3684 2 1 3800 3806 3841 3706 3840 3829 3828 1299 ICV_13 $T=642320 1041720 0 180 $X=637980 $Y=1036300
X4873 4509 4505 2 1 4438 4413 4555 4543 4550 724 4487 1299 ICV_13 $T=766940 1011480 0 180 $X=762600 $Y=1006060
X4874 4450 4446 2 1 4449 4432 4555 4543 4564 4425 4424 1299 ICV_13 $T=768800 1001400 1 180 $X=764460 $Y=1001020
X4875 4529 4539 2 1 4472 4533 4576 4540 4598 4484 4506 1299 ICV_13 $T=773140 961080 0 180 $X=768800 $Y=955660
X4876 755 748 2 1 4508 4545 4579 758 4608 757 4460 1299 ICV_13 $T=774380 910680 1 180 $X=770040 $Y=910300
X4877 5049 851 2 1 5008 5018 4959 4995 5066 879 5048 1299 ICV_13 $T=848780 920760 0 180 $X=844440 $Y=915340
X4878 5089 880 2 1 884 868 883 886 893 890 887 1299 ICV_13 $T=855600 1082040 1 180 $X=851260 $Y=1081660
X4879 5190 5138 2 1 5165 4703 4997 4992 5220 5175 5193 1299 ICV_13 $T=872340 951000 1 180 $X=868000 $Y=950620
X4880 5230 5245 2 1 5188 4934 5248 5214 5210 5244 5199 1299 ICV_13 $T=879780 1061880 1 180 $X=875440 $Y=1061500
X4881 5444 5442 2 1 5398 970 5465 5453 5456 5443 965 1299 ICV_13 $T=918840 1041720 1 180 $X=914500 $Y=1041340
X4882 5514 5442 2 1 5493 5395 5465 5453 5530 5515 977 1299 ICV_13 $T=931240 1041720 1 180 $X=926900 $Y=1041340
X4883 5640 5627 2 1 5583 5575 5655 5644 5651 1027 5623 1299 ICV_13 $T=948600 1061880 1 180 $X=944260 $Y=1061500
X4884 5728 5603 2 1 5686 5498 5687 5636 5742 5691 5724 1299 ICV_13 $T=965960 951000 1 180 $X=961620 $Y=950620
X4885 5843 1084 2 1 1082 5718 5892 5877 1093 1089 5868 1299 ICV_13 $T=996340 1082040 1 180 $X=992000 $Y=1081660
X4886 5933 1108 2 1 5863 5809 1116 1113 5952 5941 5924 1299 ICV_13 $T=1006260 1061880 1 180 $X=1001920 $Y=1061500
X4887 6117 1160 2 1 6049 1121 1168 1165 5919 6098 6079 1299 ICV_13 $T=1038500 1071960 1 180 $X=1034160 $Y=1071580
X4888 6279 6265 2 1 6264 6227 6192 6277 6292 6209 6284 1299 ICV_13 $T=1072600 1031640 1 180 $X=1068260 $Y=1031260
X4889 6269 6265 2 1 6272 1176 6192 6277 6305 6281 6243 1299 ICV_13 $T=1073840 1021560 0 180 $X=1069500 $Y=1016140
X4890 6368 1234 2 1 6337 6330 1243 6378 6379 6373 6291 1299 ICV_13 $T=1091200 1021560 0 180 $X=1086860 $Y=1016140
X4891 236 1 2 2614 2571 2588 1299 ICV_14 $T=412920 1071960 1 0 $X=412920 $Y=1066540
X4892 3391 1 2 3559 3524 3526 1299 ICV_14 $T=585280 1041720 0 0 $X=585280 $Y=1041340
X4893 3846 1 2 3927 3884 3877 1299 ICV_14 $T=654100 1001400 1 0 $X=654100 $Y=995980
X4894 3854 1 2 4114 4076 4094 1299 ICV_14 $T=684480 920760 1 0 $X=684480 $Y=915340
X4895 4058 1 2 4153 4115 4136 1299 ICV_14 $T=691300 930840 0 0 $X=691300 $Y=930460
X4896 4148 1 2 4161 4040 4073 1299 ICV_14 $T=692540 1031640 0 0 $X=692540 $Y=1031260
X4897 643 1 2 4231 657 4215 1299 ICV_14 $T=704320 1082040 0 0 $X=704320 $Y=1081660
X4898 4343 1 2 4423 4356 4391 1299 ICV_14 $T=737800 1001400 0 0 $X=737800 $Y=1001020
X4899 4446 1 2 4461 4424 4447 1299 ICV_14 $T=745860 971160 1 0 $X=745860 $Y=965740
X4900 4540 1 2 4543 4514 4534 1299 ICV_14 $T=762600 981240 1 0 $X=762600 $Y=975820
X4901 4501 1 2 4493 4502 4535 1299 ICV_14 $T=766320 1051800 1 0 $X=766320 $Y=1046380
X4902 4541 1 2 4592 4612 4641 1299 ICV_14 $T=783060 1011480 1 0 $X=783060 $Y=1006060
X4903 4922 1 2 4971 4874 4930 1299 ICV_14 $T=828320 930840 0 0 $X=828320 $Y=930460
X4904 868 1 2 975 5412 5434 1299 ICV_14 $T=910780 1082040 0 0 $X=910780 $Y=1081660
X4905 5508 1 2 5452 5488 5511 1299 ICV_14 $T=924420 1031640 1 0 $X=924420 $Y=1026220
X4906 5497 1 2 5528 5638 5662 1299 ICV_14 $T=949220 1001400 1 0 $X=949220 $Y=995980
X4907 6093 1 2 6144 6032 6095 1299 ICV_14 $T=1050900 1021560 0 0 $X=1050900 $Y=1021180
X4908 6162 1 2 6259 6224 6262 1299 ICV_14 $T=1066400 981240 1 0 $X=1066400 $Y=975820
X4909 6246 1 2 6271 6237 6218 1299 ICV_14 $T=1070740 900600 0 0 $X=1070740 $Y=900220
X4910 6348 1 2 1241 1232 1236 1299 ICV_14 $T=1086240 900600 0 0 $X=1086240 $Y=900220
X4911 226 1 2 230 2462 185 223 2502 1299 ICV_15 $T=394320 1082040 0 0 $X=394320 $Y=1081660
X4912 2797 1 2 2820 2732 253 2753 2774 1299 ICV_15 $T=438340 951000 1 0 $X=438340 $Y=945580
X4913 315 1 2 319 2881 252 309 298 1299 ICV_15 $T=472440 1082040 0 0 $X=472440 $Y=1081660
X4914 2975 1 2 2969 2936 253 2875 2965 1299 ICV_15 $T=475540 930840 0 0 $X=475540 $Y=930460
X4915 3008 1 2 3040 3103 252 3071 3153 1299 ICV_15 $T=506540 1051800 1 0 $X=506540 $Y=1046380
X4916 3183 1 2 3162 3130 253 3134 3183 1299 ICV_15 $T=510880 940920 1 0 $X=510880 $Y=935500
X4917 364 1 2 368 3136 252 360 3160 1299 ICV_15 $T=512120 1082040 0 0 $X=512120 $Y=1081660
X4918 377 1 2 389 3196 253 3228 2365 1299 ICV_15 $T=523280 930840 1 0 $X=523280 $Y=925420
X4919 3329 1 2 3363 3274 380 3294 3299 1299 ICV_15 $T=538160 930840 0 0 $X=538160 $Y=930460
X4920 3416 1 2 3438 3346 2637 3391 3410 1299 ICV_15 $T=550560 1051800 1 0 $X=550560 $Y=1046380
X4921 3410 1 2 3411 3360 399 3356 3357 1299 ICV_15 $T=552420 1071960 1 0 $X=552420 $Y=1066540
X4922 3514 1 2 3504 3465 380 3407 3514 1299 ICV_15 $T=571640 951000 0 0 $X=571640 $Y=950620
X4923 3865 1 2 3864 3810 380 3821 3573 1299 ICV_15 $T=639220 940920 1 0 $X=639220 $Y=935500
X4924 4092 1 2 4090 4035 599 4019 632 1299 ICV_15 $T=677660 1061880 0 0 $X=677660 $Y=1061500
X4925 827 1 2 839 4773 799 804 4805 1299 ICV_15 $T=801040 1082040 0 0 $X=801040 $Y=1081660
X4926 5074 1 2 5056 5019 4870 5067 879 1299 ICV_15 $T=845680 930840 0 0 $X=845680 $Y=930460
X4927 5236 1 2 5229 5178 869 915 5236 1299 ICV_15 $T=869860 910680 1 0 $X=869860 $Y=905260
X4928 5504 1 2 5540 5467 5328 5451 5529 1299 ICV_15 $T=921320 1021560 0 0 $X=921320 $Y=1021180
X4929 5501 1 2 5543 5481 946 5560 5407 1299 ICV_15 $T=929380 1061880 1 0 $X=929380 $Y=1056460
X4930 5769 1 2 5788 5738 5328 5717 5769 1299 ICV_15 $T=966580 1021560 1 0 $X=966580 $Y=1016140
X4931 5472 1 2 5470 6054 1115 6018 1132 1299 ICV_15 $T=1027960 920760 0 0 $X=1027960 $Y=920380
X4932 6149 1 2 6112 6087 6041 6029 6149 1299 ICV_15 $T=1034160 961080 0 0 $X=1034160 $Y=960700
X4933 6210 1 2 6204 6161 6041 6126 6171 1299 ICV_15 $T=1047800 981240 1 0 $X=1047800 $Y=975820
X4934 6228 1 2 6234 6176 1149 1198 6228 1299 ICV_15 $T=1052140 1061880 1 0 $X=1052140 $Y=1056460
X4935 6244 1 2 6214 6245 6041 6162 1211 1299 ICV_15 $T=1063920 951000 1 0 $X=1063920 $Y=945580
X4936 6350 1 2 6334 6307 1115 6312 1233 1299 ICV_15 $T=1078800 930840 0 0 $X=1078800 $Y=930460
X4937 6395 1 2 6423 6340 1149 1235 6386 1299 ICV_15 $T=1085000 1082040 1 0 $X=1085000 $Y=1076620
X4938 87 2 49 1 87 1920 1299 ICV_16 $T=308140 940920 0 0 $X=308140 $Y=940540
X4939 1920 2 1615 1 1920 135 1299 ICV_16 $T=331700 940920 0 0 $X=331700 $Y=940540
X4940 3157 2 3253 1 3253 3144 1299 ICV_16 $T=533820 1001400 1 0 $X=533820 $Y=995980
X4941 621 2 4060 1 4060 4191 1299 ICV_16 $T=701840 1021560 1 0 $X=701840 $Y=1016140
X4942 4524 2 739 1 621 4524 1299 ICV_16 $T=765700 910680 1 0 $X=765700 $Y=905260
X4943 4782 2 5010 1 5010 5021 1299 ICV_16 $T=841960 991320 1 0 $X=841960 $Y=985900
X4944 5183 2 5204 1 4607 5214 1299 ICV_16 $T=873580 1031640 0 0 $X=873580 $Y=1031260
X4945 5280 2 5399 1 5280 5391 1299 ICV_16 $T=906440 940920 0 0 $X=906440 $Y=940540
X4946 5553 2 5571 1 5571 5558 1299 ICV_16 $T=938060 930840 0 0 $X=938060 $Y=930460
X4947 5505 2 5609 1 5572 5635 1299 ICV_16 $T=947360 940920 1 0 $X=947360 $Y=935500
X4948 841 2 5683 1 5683 5718 1299 ICV_16 $T=959760 1082040 0 0 $X=959760 $Y=1081660
X4949 6002 2 6004 1 5598 6014 1299 ICV_16 $T=1017420 1001400 0 0 $X=1017420 $Y=1001020
X4950 5910 2 6031 1 6031 1118 1299 ICV_16 $T=1021760 1061880 0 0 $X=1021760 $Y=1061500
X4951 1099 2 6052 1 6052 6060 1299 ICV_16 $T=1027340 981240 1 0 $X=1027340 $Y=975820
X4952 6187 2 6230 1 6230 6236 1299 ICV_16 $T=1061440 1031640 0 0 $X=1061440 $Y=1031260
X4953 6201 2 6249 1 6249 6255 1299 ICV_16 $T=1064540 991320 1 0 $X=1064540 $Y=985900
X4954 1216 2 1173 1 6261 1212 1299 ICV_16 $T=1078800 920760 1 0 $X=1078800 $Y=915340
X4955 2317 2 189 1 2290 2324 1299 ICV_17 $T=368900 981240 0 0 $X=368900 $Y=980860
X4956 2373 2 2380 1 2348 2369 1299 ICV_17 $T=376340 1031640 1 0 $X=376340 $Y=1026220
X4957 2380 2 2377 1 2383 2409 1299 ICV_17 $T=382540 1001400 0 0 $X=382540 $Y=1001020
X4958 2478 2 2507 1 2477 2499 1299 ICV_17 $T=397420 981240 1 0 $X=397420 $Y=975820
X4959 2872 2 2957 1 2920 2930 1299 ICV_17 $T=473680 1071960 1 0 $X=473680 $Y=1066540
X4960 3079 2 3316 1 3236 3247 1299 ICV_17 $T=537540 991320 1 0 $X=537540 $Y=985900
X4961 3559 2 3646 1 3611 3640 1299 ICV_17 $T=603880 1021560 0 0 $X=603880 $Y=1021180
X4962 3582 2 3711 1 3650 3686 1299 ICV_17 $T=613800 1001400 1 0 $X=613800 $Y=995980
X4963 580 2 587 1 3898 3925 1299 ICV_17 $T=656580 940920 0 0 $X=656580 $Y=940540
X4964 3904 2 4025 1 3982 4007 1299 ICV_17 $T=669600 930840 0 0 $X=669600 $Y=930460
X4965 3316 2 4134 1 4224 4267 1299 ICV_17 $T=714860 991320 1 0 $X=714860 $Y=985900
X4966 5187 2 5233 1 5192 5226 1299 ICV_17 $T=873580 1021560 1 0 $X=873580 $Y=1016140
X4967 5351 2 5354 1 5309 5348 1299 ICV_17 $T=892180 1051800 1 0 $X=892180 $Y=1046380
X4968 5804 2 5922 1 5884 5913 1299 ICV_17 $T=999440 1021560 1 0 $X=999440 $Y=1016140
X4969 5922 2 5975 1 5974 6011 1299 ICV_17 $T=1014320 1021560 0 0 $X=1014320 $Y=1021180
X4970 6200 2 6201 1 6171 6193 1299 ICV_17 $T=1052760 961080 0 0 $X=1052760 $Y=960700
X4971 2469 2298 1 2 INV6CK $T=396800 1041720 0 180 $X=391220 $Y=1036300
X4972 250 2469 1 2 INV6CK $T=432760 1031640 0 180 $X=427180 $Y=1026220
X4973 247 250 1 2 INV6CK $T=430280 1011480 0 0 $X=430280 $Y=1011100
X4974 3673 576 1 2 INV6CK $T=652240 961080 0 0 $X=652240 $Y=960700
X4975 4918 5711 1 2 INV6CK $T=967200 1021560 0 0 $X=967200 $Y=1021180
X4976 4918 5964 1 2 INV6CK $T=1008120 1021560 0 0 $X=1008120 $Y=1021180
X4977 5925 1110 1104 5919 5471 1 2 AN4 $T=1007500 1082040 0 180 $X=1001300 $Y=1076620
X4978 4684 912 5228 5231 2 1 NR3H $T=876060 1031640 0 0 $X=876060 $Y=1031260
X4979 3997 5422 5494 998 2 1 NR3H $T=924420 971160 0 0 $X=924420 $Y=970780
X4980 1322 1320 1300 1 2 ND2 $T=222580 1011480 1 180 $X=220720 $Y=1011100
X4981 1321 1311 1325 1 2 ND2 $T=222580 1051800 0 0 $X=222580 $Y=1051420
X4982 1323 1355 1340 1 2 ND2 $T=228160 1011480 0 180 $X=226300 $Y=1006060
X4983 2777 2778 2515 1 2 ND2 $T=446400 1001400 0 180 $X=444540 $Y=995980
X4984 2958 2954 2730 1 2 ND2 $T=479880 940920 1 180 $X=478020 $Y=940540
X4985 4647 4644 4568 1 2 ND2 $T=783680 1051800 1 0 $X=783680 $Y=1046380
X4986 4661 4631 4639 1 2 ND2 $T=785540 1041720 0 0 $X=785540 $Y=1041340
X4987 5371 5410 5255 1 2 ND2 $T=910160 940920 0 0 $X=910160 $Y=940540
X4988 4653 4789 4797 4809 2 1 4821 OA112 $T=803520 1021560 1 0 $X=803520 $Y=1016140
X4989 4548 4799 4797 4815 2 1 4827 OA112 $T=804140 1031640 0 0 $X=804140 $Y=1031260
X4990 4602 4816 4797 4832 2 1 4841 OA112 $T=806000 1061880 1 0 $X=806000 $Y=1056460
X4991 4630 4820 4797 4837 2 1 4842 OA112 $T=806620 1011480 1 0 $X=806620 $Y=1006060
X4992 4594 4844 4797 4829 2 1 4866 OA112 $T=810340 1041720 0 0 $X=810340 $Y=1041340
X4993 5184 5112 5054 5177 2 1 5215 OA112 $T=871100 1041720 1 0 $X=871100 $Y=1036300
X4994 5250 5076 5054 5233 2 1 5294 OA112 $T=881640 1011480 0 0 $X=881640 $Y=1011100
X4995 5297 5142 5054 5318 2 1 5324 OA112 $T=887840 1011480 0 0 $X=887840 $Y=1011100
X4996 5341 5107 5054 5359 2 1 5363 OA112 $T=895280 1021560 1 0 $X=895280 $Y=1016140
X4997 5304 5077 5054 5354 2 1 5379 OA112 $T=895280 1041720 1 0 $X=895280 $Y=1036300
X4998 2469 3056 1 2 INV8CK $T=499100 1041720 0 180 $X=492280 $Y=1036300
X4999 3673 4918 1 2 INV8CK $T=827700 1001400 0 180 $X=820880 $Y=995980
X5000 4918 4687 1 2 INV8CK $T=825220 1021560 0 0 $X=825220 $Y=1021180
X5001 3673 854 1 2 INV8CK $T=827080 910680 0 0 $X=827080 $Y=910300
X5002 4897 836 1 4880 838 4877 2 OAI112HS $T=820880 910680 1 180 $X=816540 $Y=910300
X5003 4568 4591 2 4614 767 4639 1 AOI22HP $T=770660 1031640 1 0 $X=770660 $Y=1026220
X5004 4568 4699 2 4726 798 4639 1 AOI22HP $T=802900 1021560 1 180 $X=789880 $Y=1021180
X5005 4568 4634 2 4639 776 4663 1 AOI22H $T=779960 1031640 0 0 $X=779960 $Y=1031260
X5006 4568 4680 2 4639 777 4650 1 AOI22H $T=791120 1031640 0 180 $X=783680 $Y=1026220
X5007 4568 4700 2 4688 786 4639 1 AOI22H $T=794840 1051800 0 180 $X=787400 $Y=1046380
X5008 4684 4614 3870 791 1 2 ND3P $T=787400 1031640 0 0 $X=787400 $Y=1031260
X5009 3713 2 3517 1 3736 NR2P $T=624340 1051800 1 180 $X=620620 $Y=1051420
X5010 3859 2 3395 1 3870 NR2P $T=652240 1051800 1 180 $X=648520 $Y=1051420
X5011 3875 2 569 1 3881 NR2P $T=650380 1051800 1 0 $X=650380 $Y=1046380
X5012 1953 120 85 2 121 1 124 AN4B1S $T=321780 1082040 0 0 $X=321780 $Y=1081660
X5013 3242 3234 3205 2 2669 1 3224 AN4B1S $T=533820 1001400 0 180 $X=529480 $Y=995980
X5014 3289 3282 3239 2 3049 1 3272 AN4B1S $T=542500 971160 1 180 $X=538160 $Y=970780
X5015 3319 3310 3237 2 3039 1 3295 AN4B1S $T=546840 951000 1 180 $X=542500 $Y=950620
X5016 3326 3331 3173 2 2610 1 3325 AN4B1S $T=549940 1001400 0 180 $X=545600 $Y=995980
X5017 3384 3393 3238 2 2839 1 3406 AN4B1S $T=558000 951000 1 0 $X=558000 $Y=945580
X5018 3426 3430 3244 2 2596 1 3449 AN4B1S $T=564200 991320 1 0 $X=564200 $Y=985900
X5019 3455 3459 3341 2 2808 1 3470 AN4B1S $T=569780 951000 1 0 $X=569780 $Y=945580
X5020 3482 3476 3216 2 2796 1 3463 AN4B1S $T=575980 971160 1 180 $X=571640 $Y=970780
X5021 3480 3484 3226 2 2982 1 3471 AN4B1S $T=577840 961080 0 180 $X=573500 $Y=955660
X5022 3503 3498 3418 2 453 1 454 AN4B1S $T=582180 900600 1 180 $X=577840 $Y=900220
X5023 3477 3497 3227 2 2886 1 3509 AN4B1S $T=578460 991320 1 0 $X=578460 $Y=985900
X5024 3528 3518 3456 2 2928 1 461 AN4B1S $T=585900 920760 0 180 $X=581560 $Y=915340
X5025 3564 3541 3381 2 2932 1 480 AN4B1S $T=594580 920760 1 180 $X=590240 $Y=920380
X5026 312 1 2 2540 BUF3CK $T=483600 940920 0 0 $X=483600 $Y=940540
X5027 1337 2 1376 1318 1307 1 1301 FA1S $T=231880 910680 0 180 $X=220100 $Y=905260
X5028 7 2 13 15 1337 1 1305 FA1S $T=232500 900600 1 180 $X=220720 $Y=900220
X5029 8 2 1381 12 1362 1 1303 FA1S $T=232500 910680 1 180 $X=220720 $Y=910300
X5030 9 2 1404 1356 1370 1 1312 FA1S $T=233120 930840 0 180 $X=221340 $Y=925420
X5031 1351 2 1328 1343 1371 1 1313 FA1S $T=233120 940920 0 180 $X=221340 $Y=935500
X5032 6 2 1329 1305 1349 1 1330 FA1S $T=221340 951000 1 0 $X=221340 $Y=945580
X5033 1349 2 1352 1344 1372 1 1314 FA1S $T=233120 961080 0 180 $X=221340 $Y=955660
X5034 1335 2 1354 1392 1331 1 1302 FA1S $T=233120 1031640 1 180 $X=221340 $Y=1031260
X5035 1336 2 1359 1327 1384 1 1394 FA1S $T=222580 1061880 0 0 $X=222580 $Y=1061500
X5036 1365 2 1421 1435 1411 1 1347 FA1S $T=238700 1051800 0 180 $X=226920 $Y=1046380
X5037 1370 2 1379 1458 1414 1 1357 FA1S $T=240560 930840 1 180 $X=228780 $Y=930460
X5038 1372 2 1390 1426 1415 1 1348 FA1S $T=240560 951000 1 180 $X=228780 $Y=950620
X5039 1381 2 1457 1424 1428 1 1363 FA1S $T=241180 920760 0 180 $X=229400 $Y=915340
X5040 1371 2 1382 1425 1407 1 1366 FA1S $T=241800 940920 1 180 $X=230020 $Y=940540
X5041 1411 2 1393 1441 1430 1 1368 FA1S $T=241800 1051800 1 180 $X=230020 $Y=1051420
X5042 1420 2 1396 1419 1432 1 1373 FA1S $T=242420 961080 1 180 $X=230640 $Y=960700
X5043 1427 2 1459 1373 1437 1 1377 FA1S $T=243040 981240 0 180 $X=231260 $Y=975820
X5044 1307 2 1465 1456 1436 1 1390 FA1S $T=245520 910680 1 180 $X=233740 $Y=910300
X5045 19 2 21 1466 16 1 1385 FA1S $T=246760 900600 1 180 $X=234980 $Y=900220
X5046 1353 2 1420 1398 1427 1 1433 FA1S $T=235600 971160 0 0 $X=235600 $Y=970780
X5047 1375 2 1498 1422 1462 1 1399 FA1S $T=247380 1061880 0 180 $X=235600 $Y=1056460
X5048 20 2 1454 17 1418 1 1409 FA1S $T=248000 910680 0 180 $X=236220 $Y=905260
X5049 1443 2 1406 1399 1479 1 1485 FA1S $T=236220 1071960 0 0 $X=236220 $Y=1071580
X5050 1444 2 1484 1492 1468 1 1382 FA1S $T=248620 930840 0 180 $X=236840 $Y=925420
X5051 1407 2 1445 1481 1473 1 1419 FA1S $T=249240 940920 0 180 $X=237460 $Y=935500
X5052 1467 2 1448 1488 1482 1 1422 FA1S $T=249860 1041720 0 180 $X=238080 $Y=1036300
X5053 1436 2 1487 1526 1475 1 1431 FA1S $T=250480 951000 0 180 $X=238700 $Y=945580
X5054 1464 2 1506 1524 1483 1 1354 FA1S $T=251100 1021560 0 180 $X=239320 $Y=1016140
X5055 1384 2 1505 1412 1539 1 1518 FA1S $T=240560 1061880 0 0 $X=240560 $Y=1061500
X5056 1415 2 1431 1455 1503 1 1440 FA1S $T=252960 961080 0 180 $X=241180 $Y=955660
X5057 1492 2 1527 1519 1508 1 1450 FA1S $T=254200 920760 1 180 $X=242420 $Y=920380
X5058 1475 2 1551 1530 1516 1 1460 FA1S $T=255440 951000 1 180 $X=243660 $Y=950620
X5059 1459 2 1521 1476 1532 1 1469 FA1S $T=256680 981240 0 180 $X=244900 $Y=975820
X5060 1498 2 1563 1535 1525 1 1470 FA1S $T=256680 1051800 1 180 $X=244900 $Y=1051420
X5061 1414 2 1557 1493 1543 1 1471 FA1S $T=258540 930840 1 180 $X=246760 $Y=930460
X5062 1503 2 1480 1460 1562 1 1517 FA1S $T=246760 971160 1 0 $X=246760 $Y=965740
X5063 1437 2 1565 1469 1594 1 1577 FA1S $T=249860 981240 0 0 $X=249860 $Y=980860
X5064 1462 2 1580 1547 1556 1 1497 FA1S $T=261640 1061880 0 180 $X=249860 $Y=1056460
X5065 1362 2 1583 1573 1564 1 1484 FA1S $T=262880 930840 0 180 $X=251100 $Y=925420
X5066 1479 2 1470 1497 1598 1 1561 FA1S $T=251100 1071960 0 0 $X=251100 $Y=1071580
X5067 1532 2 1571 1536 1587 1 1624 FA1S $T=252960 971160 0 0 $X=252960 $Y=970780
X5068 1454 2 35 1600 1593 1 1486 FA1S $T=265980 910680 0 180 $X=254200 $Y=905260
X5069 1515 2 1599 1502 1603 1 1625 FA1S $T=254200 1082040 0 0 $X=254200 $Y=1081660
X5070 1418 2 1621 1641 1588 1 1529 FA1S $T=266600 910680 1 180 $X=254820 $Y=910300
X5071 1432 2 1622 1575 1590 1 1521 FA1S $T=266600 951000 0 180 $X=254820 $Y=945580
X5072 1531 2 1633 1552 1597 1 1536 FA1S $T=267220 961080 1 180 $X=255440 $Y=960700
X5073 1594 2 1559 1637 1611 1 1546 FA1S $T=268460 991320 0 180 $X=256680 $Y=985900
X5074 1598 2 1635 1616 1606 1 1549 FA1S $T=268460 1061880 1 180 $X=256680 $Y=1061500
X5075 42 2 1631 52 45 1 36 FA1S $T=269080 900600 1 180 $X=257300 $Y=900220
X5076 1565 2 1651 1624 1634 1 1559 FA1S $T=271560 981240 0 180 $X=259780 $Y=975820
X5077 1603 2 1569 1518 1693 1 1658 FA1S $T=259780 1082040 1 0 $X=259780 $Y=1076620
X5078 1473 2 1655 1670 1614 1 1575 FA1S $T=272800 930840 1 180 $X=261020 $Y=930460
X5079 1562 2 1683 1663 1628 1 1581 FA1S $T=275280 971160 0 180 $X=263500 $Y=965740
X5080 1637 2 1607 1668 1699 1 1691 FA1S $T=264740 981240 0 0 $X=264740 $Y=980860
X5081 1587 2 1709 1623 1675 1 1607 FA1S $T=279000 971160 1 180 $X=267220 $Y=970780
X5082 1611 2 1704 1691 1680 1 1629 FA1S $T=280240 1001400 0 180 $X=268460 $Y=995980
X5083 58 2 1703 1714 1694 1 1641 FA1S $T=281480 910680 1 180 $X=269700 $Y=910300
X5084 1539 2 1708 1705 1701 1 1645 FA1S $T=282100 1061880 1 180 $X=270320 $Y=1061500
X5085 1693 2 1645 1712 1710 1 1649 FA1S $T=282720 1071960 0 180 $X=270940 $Y=1066540
X5086 1680 2 1660 1706 1775 1 1740 FA1S $T=271560 991320 1 0 $X=271560 $Y=985900
X5087 1468 2 1741 1732 1721 1 1481 FA1S $T=285820 930840 1 180 $X=274040 $Y=930460
X5088 1590 2 1739 1753 1722 1 1634 FA1S $T=285820 951000 0 180 $X=274040 $Y=945580
X5089 1668 2 1696 1679 1728 1 1660 FA1S $T=285820 981240 0 180 $X=274040 $Y=975820
X5090 1653 2 1667 1649 1766 1 1752 FA1S $T=274660 1071960 0 0 $X=274660 $Y=1071580
X5091 1583 2 1748 1738 1743 1 1508 FA1S $T=288300 920760 0 180 $X=276520 $Y=915340
X5092 1631 2 1770 1788 1756 1 1466 FA1S $T=291400 900600 1 180 $X=279620 $Y=900220
X5093 1699 2 1797 1713 1755 1 1706 FA1S $T=291400 981240 1 180 $X=279620 $Y=980860
X5094 1721 2 1795 1798 1750 1 1655 FA1S $T=292640 930840 0 180 $X=280860 $Y=925420
X5095 1675 2 1786 1715 1747 1 1713 FA1S $T=292640 971160 0 180 $X=280860 $Y=965740
X5096 1756 2 65 1729 1725 1 1621 FA1S $T=293260 910680 0 180 $X=281480 $Y=905260
X5097 1651 2 1794 1759 1673 1 1704 FA1S $T=293880 971160 1 180 $X=282100 $Y=970780
X5098 1606 2 1761 1792 1801 1 1815 FA1S $T=283960 1061880 0 0 $X=283960 $Y=1061500
X5099 1766 2 1719 1809 1838 1 1825 FA1S $T=285200 1071960 1 0 $X=285200 $Y=1066540
X5100 1710 2 1783 1751 1773 1 1837 FA1S $T=285820 1061880 1 0 $X=285820 $Y=1056460
X5101 1775 2 1760 1802 1830 1 1834 FA1S $T=286440 991320 0 0 $X=286440 $Y=990940
X5102 1564 2 1840 1803 1805 1 1732 FA1S $T=300700 920760 1 180 $X=288920 $Y=920380
X5103 1526 2 1852 1781 1833 1 1731 FA1S $T=301320 951000 0 180 $X=289540 $Y=945580
X5104 1755 2 1698 1860 1843 1 1760 FA1S $T=301320 981240 0 180 $X=289540 $Y=975820
X5105 1788 2 78 1864 1839 1 1600 FA1S $T=304420 900600 1 180 $X=292640 $Y=900220
X5106 1830 2 1867 1727 1884 1 1878 FA1S $T=294500 981240 0 0 $X=294500 $Y=980860
X5107 1665 2 1886 1817 1949 1 1908 FA1S $T=297600 1082040 1 0 $X=297600 $Y=1076620
X5108 1588 2 1925 1919 1909 1 1527 FA1S $T=312480 910680 1 180 $X=300700 $Y=910300
X5109 1890 2 1841 1851 1882 1 1945 FA1S $T=301320 1061880 1 0 $X=301320 $Y=1056460
X5110 1886 2 1857 1846 1890 1 1934 FA1S $T=301320 1071960 1 0 $X=301320 $Y=1066540
X5111 1843 2 1861 1819 1875 1 1867 FA1S $T=302560 971160 0 0 $X=302560 $Y=970780
X5112 1838 2 1899 1891 1951 1 1940 FA1S $T=309380 1061880 0 0 $X=309380 $Y=1061500
X5113 1949 2 1979 1934 1981 1 1999 FA1S $T=311860 1071960 0 0 $X=311860 $Y=1071580
X5114 1770 2 103 1942 109 1 1593 FA1S $T=312480 900600 0 0 $X=312480 $Y=900220
X5115 1971 2 1956 1885 1954 1 2064 FA1S $T=315580 1061880 1 0 $X=315580 $Y=1056460
X5116 1981 2 1945 1946 1971 1 2027 FA1S $T=318060 1071960 1 0 $X=318060 $Y=1066540
X5117 2057 2 2032 2103 2068 1 2005 FA1S $T=337900 991320 1 180 $X=326120 $Y=990940
X5118 2063 2 2072 2094 2073 1 2010 FA1S $T=338520 981240 0 180 $X=326740 $Y=975820
X5119 2069 2 2057 2087 2077 1 1964 FA1S $T=339140 1001400 0 180 $X=327360 $Y=995980
X5120 2074 2 1879 2017 2130 1 2114 FA1S $T=330460 1041720 1 0 $X=330460 $Y=1036300
X5121 2026 2 2074 2012 2064 1 2119 FA1S $T=330460 1051800 0 0 $X=330460 $Y=1051420
X5122 2089 2 2133 2102 2080 1 2043 FA1S $T=342860 981240 1 180 $X=331080 $Y=980860
X5123 2077 2 2050 2063 2089 1 2103 FA1S $T=331080 991320 1 0 $X=331080 $Y=985900
X5124 2078 2 2036 2114 2049 1 2122 FA1S $T=331080 1041720 0 0 $X=331080 $Y=1041340
X5125 2079 2 2078 2119 2107 1 2037 FA1S $T=343480 1051800 0 180 $X=331700 $Y=1046380
X5126 2106 2 2143 1955 2022 1 2102 FA1S $T=335420 961080 0 0 $X=335420 $Y=960700
X5127 2127 2 2168 2132 2106 1 2050 FA1S $T=347820 971160 1 180 $X=336040 $Y=970780
X5128 2126 2 2004 2116 2124 1 2172 FA1S $T=338520 951000 0 0 $X=338520 $Y=950620
X5129 154 2 2120 143 2051 1 2192 FA1S $T=339760 920760 1 0 $X=339760 $Y=915340
X5130 2068 2 2010 2043 2166 1 2179 FA1S $T=340380 991320 0 0 $X=340380 $Y=990940
X5131 2147 2 2169 152 149 1 2195 FA1S $T=341000 910680 1 0 $X=341000 $Y=905260
X5132 2148 2 2141 2131 2113 1 2187 FA1S $T=341000 930840 0 0 $X=341000 $Y=930460
X5133 2107 2 2214 2122 2193 1 2139 FA1S $T=356500 1031640 1 180 $X=344720 $Y=1031260
X5134 2166 2 2138 2152 2181 1 2190 FA1S $T=345340 991320 1 0 $X=345340 $Y=985900
X5135 2170 2 170 2099 2147 1 2226 FA1S $T=345960 910680 0 0 $X=345960 $Y=910300
X5136 2181 2 2162 2048 2173 1 2167 FA1S $T=347200 981240 0 0 $X=347200 $Y=980860
X5137 2207 2 2188 2238 2067 1 2162 FA1S $T=360220 961080 1 180 $X=348440 $Y=960700
X5138 2080 2 2062 2223 2207 1 2138 FA1S $T=360840 971160 0 180 $X=349060 $Y=965740
X5139 2199 2 167 165 2206 1 2225 FA1S $T=349680 920760 0 0 $X=349680 $Y=920380
X5140 2206 2 2148 163 2235 1 2246 FA1S $T=350300 930840 1 0 $X=350300 $Y=925420
X5141 2230 2 2249 2247 1987 1 2032 FA1S $T=363940 971160 1 180 $X=352160 $Y=970780
X5142 2221 2 176 2195 2101 1 2268 FA1S $T=352780 900600 0 0 $X=352780 $Y=900220
X5143 2232 2 2218 2202 2201 1 2283 FA1S $T=354640 1001400 0 0 $X=354640 $Y=1001020
X5144 2235 2 2060 2259 2286 1 2289 FA1S $T=355260 930840 0 0 $X=355260 $Y=930460
X5145 2214 2 2211 2178 2088 1 2291 FA1S $T=357740 1041720 1 0 $X=357740 $Y=1036300
X5146 180 2 2221 2226 179 1 2308 FA1S $T=360220 910680 0 0 $X=360220 $Y=910300
X5147 181 2 2237 2245 2321 1 2335 FA1S $T=360220 920760 1 0 $X=360220 $Y=915340
X5148 2281 2 2230 2301 2293 1 2087 FA1S $T=372000 991320 0 180 $X=360220 $Y=985900
X5149 2288 2 2281 2310 2069 1 2156 FA1S $T=373240 991320 1 180 $X=361460 $Y=990940
X5150 2273 2 2255 2312 2127 1 2301 FA1S $T=362080 981240 1 0 $X=362080 $Y=975820
X5151 2270 2 2239 2224 2232 1 2306 FA1S $T=362080 1021560 0 0 $X=362080 $Y=1021180
X5152 2279 2 2125 2253 2142 1 2312 FA1S $T=362700 961080 0 0 $X=362700 $Y=960700
X5153 2280 2 2282 2013 1967 1 2266 FA1S $T=362700 971160 1 0 $X=362700 $Y=965740
X5154 2286 2 2252 2269 2299 1 2337 FA1S $T=363940 930840 1 0 $X=363940 $Y=925420
X5155 2193 2 2244 2291 2270 1 2297 FA1S $T=363940 1031640 1 0 $X=363940 $Y=1026220
X5156 2342 2 2320 2314 2309 1 2293 FA1S $T=371380 961080 1 0 $X=371380 $Y=955660
X5157 2343 2 2338 2172 2280 1 2376 FA1S $T=371380 971160 0 0 $X=371380 $Y=970780
X5158 2259 2 2372 2315 2326 1 2388 FA1S $T=372000 910680 0 0 $X=372000 $Y=910300
X5159 2368 2 2395 2386 2353 1 2331 FA1S $T=385640 951000 1 180 $X=373860 $Y=950620
X5160 2389 2 2367 2405 2288 1 1844 FA1S $T=388120 991320 0 180 $X=376340 $Y=985900
X5161 2367 2 2354 2345 2273 1 2310 FA1S $T=376960 981240 0 0 $X=376960 $Y=980860
X5162 2397 2 2364 2404 2342 1 2354 FA1S $T=389360 961080 1 180 $X=377580 $Y=960700
X5163 2396 2 2039 2171 2399 1 2449 FA1S $T=380060 940920 0 0 $X=380060 $Y=940540
X5164 2412 2 2393 2427 2343 1 2401 FA1S $T=383160 971160 1 0 $X=383160 $Y=965740
X5165 2421 2 2375 2447 2350 1 2426 FA1S $T=385020 920760 0 0 $X=385020 $Y=920380
X5166 210 2 2363 2341 2357 1 2472 FA1S $T=385640 910680 1 0 $X=385640 $Y=905260
X5167 2451 2 2487 2368 2126 1 2393 FA1S $T=397420 961080 0 180 $X=385640 $Y=955660
X5168 2430 2 2425 2337 2421 1 2476 FA1S $T=386260 930840 1 0 $X=386260 $Y=925420
X5169 2456 2 2426 2471 2033 1 2404 FA1S $T=398040 951000 0 180 $X=386260 $Y=945580
X5170 2439 2 2407 2418 2397 1 2405 FA1S $T=386880 971160 0 0 $X=386880 $Y=970780
X5171 2464 2 2484 2476 2456 1 2418 FA1S $T=399900 951000 1 180 $X=388120 $Y=950620
X5172 2478 2 2439 2491 2389 1 2264 FA1S $T=402380 981240 1 180 $X=390600 $Y=980860
X5173 219 2 217 2366 2473 1 2530 FA1S $T=393700 910680 0 0 $X=393700 $Y=910300
X5174 2506 2 2525 2479 2412 1 2468 FA1S $T=407960 961080 1 180 $X=396180 $Y=960700
X5175 2504 2 2530 2472 2518 1 2557 FA1S $T=398660 920760 1 0 $X=398660 $Y=915340
X5176 2505 2 2289 2538 2430 1 2559 FA1S $T=398660 930840 0 0 $X=398660 $Y=930460
X5177 2538 2 2572 2083 2388 1 2432 FA1S $T=411680 920760 1 180 $X=399900 $Y=920380
X5178 2518 2 220 2485 222 1 2572 FA1S $T=400520 910680 1 0 $X=400520 $Y=905260
X5179 2544 2 2559 2576 2464 1 2497 FA1S $T=412920 951000 0 180 $X=401140 $Y=945580
X5180 2550 2 2507 2578 2506 1 1782 FA1S $T=414160 961080 0 180 $X=402380 $Y=955660
X5181 2547 2 2196 2537 2396 1 2593 FA1S $T=404240 940920 0 0 $X=404240 $Y=940540
X5182 2580 2 2144 238 2591 1 2542 FA1S $T=419120 910680 1 180 $X=407340 $Y=910300
X5183 2321 2 2568 2403 2547 1 2583 FA1S $T=408580 940920 1 0 $X=408580 $Y=935500
X5184 2592 2 2577 2562 2451 1 2525 FA1S $T=411060 930840 1 0 $X=411060 $Y=925420
X5185 2604 2 2580 2192 2504 1 2640 FA1S $T=412920 920760 0 0 $X=412920 $Y=920380
X5186 237 2 234 235 2475 1 2591 FA1S $T=414780 900600 0 0 $X=414780 $Y=900220
X5187 2609 2 2627 2602 2544 1 2590 FA1S $T=416020 951000 0 0 $X=416020 $Y=950620
X5188 2417 2 245 2654 2604 1 2678 FA1S $T=419740 920760 1 0 $X=419740 $Y=915340
X5189 2654 2 244 246 2268 1 2664 FA1S $T=420980 910680 0 0 $X=420980 $Y=910300
X5190 2665 2 2335 2671 2684 1 2632 FA1S $T=432760 930840 1 180 $X=420980 $Y=930460
X5191 2661 2 2616 2632 2550 1 1528 FA1S $T=421600 940920 0 0 $X=421600 $Y=940540
X5192 2684 2 2655 2646 2592 1 2636 FA1S $T=426560 930840 1 0 $X=426560 $Y=925420
X5193 1994 1992 2013 2 1 XNR2HS $T=323640 971160 0 0 $X=323640 $Y=970780
X5194 2025 2029 2088 2 1 XNR2HS $T=333560 1031640 1 0 $X=333560 $Y=1026220
X5195 2661 2665 243 2 1 XNR2HS $T=428420 940920 0 180 $X=422840 $Y=935500
X5196 1650 1647 1642 1 2 1551 OA12 $T=272800 940920 1 180 $X=269080 $Y=940540
X5197 1711 1692 1687 1 2 1505 OA12 $T=279620 1031640 0 180 $X=275900 $Y=1026220
X5198 1684 1686 1688 1 2 1708 OA12 $T=275900 1041720 0 0 $X=275900 $Y=1041340
X5199 1858 1859 1889 1 2 1543 OA12 $T=308140 930840 0 180 $X=304420 $Y=925420
X5200 91 85 88 1 2 1793 OA12 $T=310620 1082040 1 180 $X=306900 $Y=1081660
X5201 1986 1975 1960 1 2 1994 OA12 $T=322400 951000 0 0 $X=322400 $Y=950620
X5202 2002 2006 1996 1 2 2041 OA12 $T=327360 920760 1 0 $X=327360 $Y=915340
X5203 1991 2009 2031 1 2 2040 OA12 $T=327980 910680 0 0 $X=327980 $Y=910300
X5204 2045 2015 2075 1 2 2094 OA12 $T=334800 961080 1 0 $X=334800 $Y=955660
X5205 2098 141 2111 1 2 2118 OA12 $T=337900 1082040 1 0 $X=337900 $Y=1076620
X5206 2092 2065 2124 1 2 2142 OA12 $T=341620 951000 1 0 $X=341620 $Y=945580
X5207 2191 2197 2198 1 2 2224 OA12 $T=354020 1031640 1 0 $X=354020 $Y=1026220
X5208 2316 2371 2378 1 2 2399 OA12 $T=380060 930840 1 0 $X=380060 $Y=925420
X5209 2117 2489 2503 1 2 2537 OA12 $T=403620 940920 1 0 $X=403620 $Y=935500
X5210 24 1 23 24 1424 26 2 OAI22S $T=248000 900600 0 0 $X=248000 $Y=900220
X5211 1520 1 1489 1520 1458 1494 2 OAI22S $T=254820 940920 0 180 $X=251100 $Y=935500
X5212 1496 1 1534 1548 1435 1511 2 OAI22S $T=254820 1041720 0 0 $X=254820 $Y=1041340
X5213 1511 1 1548 1584 1496 1572 2 OAI22S $T=259780 1041720 1 0 $X=259780 $Y=1036300
X5214 1620 1 1627 1592 1525 1548 2 OAI22S $T=267220 1051800 1 0 $X=267220 $Y=1046380
X5215 1632 1 1619 1604 1595 1654 2 OAI22S $T=268460 920760 0 0 $X=268460 $Y=920380
X5216 1685 1 1601 1685 1679 1697 2 OAI22S $T=276520 961080 0 0 $X=276520 $Y=960700
X5217 1702 1 1576 1702 1700 56 2 OAI22S $T=281480 951000 1 180 $X=277760 $Y=950620
X5218 1718 1 1720 1718 1701 1733 2 OAI22S $T=280860 1051800 0 0 $X=280860 $Y=1051420
X5219 1876 1 1842 1900 1907 1883 2 OAI22S $T=305660 961080 0 0 $X=305660 $Y=960700
X5220 1918 1 1907 1883 1709 1900 2 OAI22S $T=311860 971160 0 180 $X=308140 $Y=965740
X5221 1929 1 1939 1625 1933 1935 2 OAI22S $T=316820 1021560 0 180 $X=313100 $Y=1016140
X5222 1937 1 1957 1953 1952 1941 2 OAI22S $T=318060 1082040 1 180 $X=314340 $Y=1081660
X5223 130 1 1957 130 1941 117 2 OAI22S $T=335420 1082040 1 180 $X=331700 $Y=1081660
X5224 2185 1 2154 2213 2168 2212 2 OAI22S $T=354020 951000 0 0 $X=354020 $Y=950620
X5225 2204 1 2149 2158 2186 150 2 OAI22S $T=358360 991320 1 180 $X=354640 $Y=990940
X5226 2212 1 2213 2229 2154 2200 2 OAI22S $T=361460 951000 1 180 $X=357740 $Y=950620
X5227 2209 1 192 2352 2323 2262 2 OAI22S $T=379440 940920 1 180 $X=375720 $Y=940540
X5228 1442 1413 1388 2 1400 1377 1 AO22 $T=238700 991320 0 180 $X=233740 $Y=985900
X5229 1395 1405 1388 2 1400 1433 1 AO22 $T=234360 1001400 1 0 $X=234360 $Y=995980
X5230 1745 1740 1618 2 1509 1723 1 AO22 $T=287060 1001400 0 180 $X=282100 $Y=995980
X5231 1791 1804 1799 2 1618 1844 1 AO22 $T=293260 1001400 1 0 $X=293260 $Y=995980
X5232 1916 1948 1799 2 1903 1964 1 AO22 $T=313720 1001400 1 0 $X=313720 $Y=995980
X5233 1966 1978 1799 2 1903 2005 1 AO22 $T=319920 1001400 1 0 $X=319920 $Y=995980
X5234 2084 2093 1935 2 1939 2037 1 AO22 $T=336660 1011480 0 0 $X=336660 $Y=1011100
X5235 2056 2053 1935 2 1939 2139 1 AO22 $T=342240 1011480 0 0 $X=342240 $Y=1011100
X5236 2254 2090 2284 2 162 2297 1 AO22 $T=365180 1011480 0 0 $X=365180 $Y=1011100
X5237 2296 2283 162 2 2284 2328 1 AO22 $T=369520 1001400 0 0 $X=369520 $Y=1001020
X5238 2347 2160 2284 2 162 2306 1 AO22 $T=375720 1011480 1 180 $X=370760 $Y=1011100
X5239 2128 2177 2204 1935 2 2317 1 2007 MUX3 $T=367040 1001400 1 0 $X=367040 $Y=995980
X5240 28 1507 1428 1 2 1493 AO12 $T=252340 910680 1 180 $X=248620 $Y=910300
X5241 1474 1523 1489 1 2 1530 AO12 $T=251720 940920 0 0 $X=251720 $Y=940540
X5242 2100 2150 2113 1 2 2171 AO12 $T=347200 940920 1 0 $X=347200 $Y=935500
X5243 144 2076 2 2120 1 2131 AOI12HS $T=341620 930840 1 0 $X=341620 $Y=925420
X5244 1324 2 1364 1315 1 AN2B1S $T=231880 1031640 0 180 $X=228780 $Y=1026220
X5245 1514 2 1510 1482 1 AN2B1S $T=252960 1041720 0 180 $X=249860 $Y=1036300
X5246 1500 2 1513 1410 1 AN2B1S $T=253580 1031640 0 180 $X=250480 $Y=1026220
X5247 1727 2 1697 1696 1 AN2B1S $T=283960 961080 1 180 $X=280860 $Y=960700
X5248 1842 2 1828 1784 1 AN2B1S $T=300080 951000 1 180 $X=296980 $Y=950620
X5249 1803 2 1828 1853 1 AN2B1S $T=298220 940920 1 0 $X=298220 $Y=935500
X5250 1983 2 1998 2025 1 AN2B1S $T=325500 1031640 1 0 $X=325500 $Y=1026220
X5251 142 2 2100 2120 1 AN2B1S $T=339760 920760 0 0 $X=339760 $Y=920380
X5252 1325 1321 1 1311 2 1300 OAI12HS $T=224440 1051800 0 180 $X=220720 $Y=1046380
X5253 1300 1322 1 1320 2 1340 OAI12HS $T=222580 1011480 0 0 $X=222580 $Y=1011100
X5254 1340 1323 1 1355 2 1380 OAI12HS $T=228780 1011480 1 0 $X=228780 $Y=1006060
X5255 1439 1443 1 1423 2 1325 OAI12HS $T=239940 1082040 0 180 $X=236220 $Y=1076620
X5256 1592 1602 1 1578 2 1421 OAI12HS $T=263500 1041720 1 180 $X=259780 $Y=1041340
X5257 1504 1579 1 1568 2 1556 OAI12HS $T=263500 1051800 1 180 $X=259780 $Y=1051420
X5258 1730 1757 1 1765 2 1722 OAI12HS $T=287060 951000 0 0 $X=287060 $Y=950620
X5259 1771 1818 1 1832 2 1741 OAI12HS $T=295120 930840 0 0 $X=295120 $Y=930460
X5260 1915 1901 1 1893 2 1882 OAI12HS $T=309380 1051800 0 180 $X=305660 $Y=1046380
X5261 2008 2021 1 2030 2 1979 OAI12HS $T=327360 1071960 0 0 $X=327360 $Y=1071580
X5262 1926 1827 1914 1898 2 1 1904 MAOI1 $T=312480 1041720 0 180 $X=307520 $Y=1036300
X5263 1707 40 2 1688 1674 1 OR3B2S $T=280240 1031640 1 180 $X=276520 $Y=1031260
X5264 1653 1658 1 1665 1599 1682 2 MOAI1 $T=270940 1082040 0 0 $X=270940 $Y=1081660
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 BUF1S $T=4340 0 0 0 $X=4340 $Y=-380
X1 5 6 3 2 7 8 MUX2 $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 5 6 QDFFRBN $T=2480 0 0 0 $X=2480 $Y=-380
X1 7 5 4 8 BUF1CK $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT BUF6CK I GND O VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=13 FDC=0
X0 1 2 3 4 INV1S $T=0 0 0 0 $X=0 $Y=-380
X1 5 6 4 7 8 9 2 MOAI1S $T=4960 0 1 180 $X=1240 $Y=-380
.ENDS
***************************************
.SUBCKT NR3HT O I3 I2 I1 VCC GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV4CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN3 I1 I2 I3 VCC GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2P I2 I1 O GND VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV3 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV3CK I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 5 NR2 $T=0 0 0 0 $X=0 $Y=-380
X1 6 2 7 8 5 NR2 $T=1860 0 0 0 $X=1860 $Y=-380
.ENDS
***************************************
.SUBCKT QDFFRBP D CK RB Q GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF2CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO13S B3 B2 B1 A1 GND VCC O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND2F I2 I1 VCC O GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO13 B3 B2 B1 A1 GND VCC O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN2T I1 I2 O GND VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND3HT I3 GND I2 I1 VCC O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2S I2 I1 VCC GND O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND2P I2 GND I1 O VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MOAI1H B1 B2 GND A1 O A2 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HA1 A B C GND VCC S
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2HS I1 I2 O VCC GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MUX2S B S VCC A GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MUX2P B S A O GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MAO222 B1 A1 C1 GND VCC O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR3 I2 I1 I3 VCC GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FA1 S B VCC A CI GND CO
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540
+ 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560
+ 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580
+ 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640
+ 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660
+ 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680
+ 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700
+ 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720
+ 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740
+ 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760
+ 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780
+ 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800
+ 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820
+ 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840
+ 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860
+ 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880
+ 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900
+ 901 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920
+ 921 922 923 924 925 926 927 928 929 930 931 932 933 934 935 936 937 938 939 940
+ 941 942 943 944 945 946 947 948 949 950 951 952 953 954 955 956 957 958 959 960
+ 961 962 963 964 965 966 967 968 969 970 971 972 973 974 975 976 977 978 979 980
+ 981 982 983 984 985 986 987 988 989 990 991 992 993 994 995 996 997 998 999 1000
+ 1001 1002 1003 1004 1005 1006 1007 1008 1009 1010 1011 1012 1013 1014 1015 1016 1017 1018 1019 1020
+ 1021 1022 1023 1024 1025 1026 1027 1028 1029 1030 1031 1032 1033 1034 1035 1036 1037 1038 1039 1040
+ 1041 1042 1043 1044 1045 1046 1047 1048 1049 1050 1051 1052 1053 1054 1055 1056 1057 1058 1059 1060
+ 1061 1062 1063 1064 1065 1066 1067 1068 1069 1070 1071 1072 1073 1074 1075 1076 1077 1078 1079 1080
+ 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 1093 1094 1095 1096 1097 1098 1099 1100
+ 1101 1102 1103 1104 1105 1106 1107 1108 1109 1110 1111 1112 1113 1114 1115 1116 1117 1118 1119 1120
+ 1121 1122 1123 1124 1125 1126 1127 1128 1129 1130 1131 1132 1133 1134 1135 1136 1137 1138 1139 1140
+ 1141 1142 1143 1144 1145 1146 1147 1148 1149 1150 1151 1152 1153 1154 1155 1156 1157 1158 1159 1160
+ 1161 1162 1163 1164 1165 1166 1167 1168 1169 1170 1171 1172 1173 1174 1175 1176 1177 1178 1179 1180
+ 1181 1182 1183 1184 1185 1186 1187 1188 1189 1190 1191 1192 1193 1194 1195 1196 1197 1198 1199 1200
+ 1201 1202 1203 1204 1205 1206 1207 1208 1209 1210 1211 1212 1213 1214 1215 1216 1217 1218 1219 1220
+ 1221 1222 1223 1224 1225 1226 1227 1228 1229 1230 1231 1232 1233 1234 1235 1236 1237 1238 1239 1240
+ 1241 1242 1243 1244 1245 1246 1247 1248 1249 1250 1251 1252 1253 1254 1255 1256 1257 1306
** N=6395 EP=1258 IP=33506 FDC=0
X0 1313 2 1310 1 INV1S $T=220100 890520 1 0 $X=220100 $Y=885100
X1 1336 2 1327 1 INV1S $T=224440 830040 1 180 $X=223200 $Y=829660
X2 1342 2 1330 1 INV1S $T=225680 850200 1 180 $X=224440 $Y=849820
X3 1350 2 1334 1 INV1S $T=225680 870360 1 180 $X=224440 $Y=869980
X4 1364 2 1402 1 INV1S $T=230640 860280 0 0 $X=230640 $Y=859900
X5 1403 2 17 1 INV1S $T=233740 900600 0 180 $X=232500 $Y=895180
X6 1451 2 1454 1 INV1S $T=241800 840120 0 0 $X=241800 $Y=839740
X7 33 2 1370 1 INV1S $T=244280 729240 1 180 $X=243040 $Y=728860
X8 1495 2 26 1 INV1S $T=249240 729240 0 180 $X=248000 $Y=723820
X9 1511 2 1482 1 INV1S $T=251100 840120 0 180 $X=249860 $Y=834700
X10 1504 2 1519 1 INV1S $T=252960 819960 0 0 $X=252960 $Y=819580
X11 1530 2 1534 1 INV1S $T=255440 809880 0 0 $X=255440 $Y=809500
X12 69 2 1581 1 INV1S $T=265360 749400 0 180 $X=264120 $Y=743980
X13 1452 2 1549 1 INV1S $T=266600 840120 1 0 $X=266600 $Y=834700
X14 1576 2 1616 1 INV1S $T=269080 799800 0 0 $X=269080 $Y=799420
X15 1593 2 1625 1 INV1S $T=270940 809880 0 0 $X=270940 $Y=809500
X16 58 2 76 1 INV1S $T=272800 819960 1 0 $X=272800 $Y=814540
X17 1565 2 1636 1 INV1S $T=273420 809880 0 0 $X=273420 $Y=809500
X18 62 2 78 1 INV1S $T=274660 830040 1 0 $X=274660 $Y=824620
X19 82 2 84 1 INV1S $T=275900 729240 0 0 $X=275900 $Y=728860
X20 72 2 1568 1 INV1S $T=275900 860280 0 0 $X=275900 $Y=859900
X21 1635 2 71 1 INV1S $T=276520 830040 1 0 $X=276520 $Y=824620
X22 1612 2 1685 1 INV1S $T=279620 830040 1 0 $X=279620 $Y=824620
X23 53 2 87 1 INV1S $T=280240 850200 0 0 $X=280240 $Y=849820
X24 1549 2 94 1 INV1S $T=284580 880440 1 0 $X=284580 $Y=875020
X25 1699 2 1724 1 INV1S $T=287680 809880 0 0 $X=287680 $Y=809500
X26 99 2 106 1 INV1S $T=288300 729240 1 0 $X=288300 $Y=723820
X27 1619 2 1726 1 INV1S $T=288300 819960 1 0 $X=288300 $Y=814540
X28 102 2 1738 1 INV1S $T=290780 850200 0 0 $X=290780 $Y=849820
X29 1786 2 1739 1 INV1S $T=294500 809880 0 180 $X=293260 $Y=804460
X30 108 2 1751 1 INV1S $T=295740 749400 0 180 $X=294500 $Y=743980
X31 110 2 90 1 INV1S $T=296980 729240 0 180 $X=295740 $Y=723820
X32 79 2 107 1 INV1S $T=295740 850200 1 0 $X=295740 $Y=844780
X33 81 2 110 1 INV1S $T=296980 729240 1 0 $X=296980 $Y=723820
X34 1796 2 112 1 INV1S $T=299460 890520 1 180 $X=298220 $Y=890140
X35 1794 2 1772 1 INV1S $T=300080 830040 0 180 $X=298840 $Y=824620
X36 1809 2 97 1 INV1S $T=304420 729240 0 0 $X=304420 $Y=728860
X37 1823 2 1777 1 INV1S $T=311860 840120 1 0 $X=311860 $Y=834700
X38 129 2 133 1 INV1S $T=311860 890520 0 0 $X=311860 $Y=890140
X39 1814 2 1851 1 INV1S $T=313720 819960 1 0 $X=313720 $Y=814540
X40 1857 2 1868 1 INV1S $T=316200 880440 0 180 $X=314960 $Y=875020
X41 153 2 116 1 INV1S $T=319920 900600 1 0 $X=319920 $Y=895180
X42 150 2 1888 1 INV1S $T=323640 729240 1 180 $X=322400 $Y=728860
X43 1607 2 1881 1 INV1S $T=322400 739320 0 0 $X=322400 $Y=738940
X44 157 2 1622 1 INV1S $T=323640 769560 1 180 $X=322400 $Y=769180
X45 1877 2 1913 1 INV1S $T=323020 759480 0 0 $X=323020 $Y=759100
X46 1849 2 136 1 INV1S $T=323020 890520 0 0 $X=323020 $Y=890140
X47 1599 2 1895 1 INV1S $T=324880 809880 0 0 $X=324880 $Y=809500
X48 1847 2 1930 1 INV1S $T=326120 739320 0 0 $X=326120 $Y=738940
X49 1613 2 1929 1 INV1S $T=326120 809880 1 0 $X=326120 $Y=804460
X50 132 2 1921 1 INV1S $T=327980 890520 0 180 $X=326740 $Y=885100
X51 1826 2 1975 1 INV1S $T=331700 789720 1 0 $X=331700 $Y=784300
X52 1976 2 1926 1 INV1S $T=332940 840120 1 180 $X=331700 $Y=839740
X53 1969 2 1638 1 INV1S $T=333560 799800 0 180 $X=332320 $Y=794380
X54 1882 2 1773 1 INV1S $T=333560 880440 1 180 $X=332320 $Y=880060
X55 1580 2 1978 1 INV1S $T=332940 799800 0 0 $X=332940 $Y=799420
X56 1976 2 1829 1 INV1S $T=335420 840120 0 180 $X=334180 $Y=834700
X57 1917 2 1993 1 INV1S $T=334800 789720 1 0 $X=334800 $Y=784300
X58 1997 2 1861 1 INV1S $T=336040 830040 1 180 $X=334800 $Y=829660
X59 1968 2 1994 1 INV1S $T=334800 880440 1 0 $X=334800 $Y=875020
X60 1564 2 2002 1 INV1S $T=336040 809880 0 0 $X=336040 $Y=809500
X61 2007 2 1976 1 INV1S $T=337280 840120 0 180 $X=336040 $Y=834700
X62 187 2 1885 1 INV1S $T=337900 789720 0 180 $X=336660 $Y=784300
X63 1982 2 2020 1 INV1S $T=339140 799800 0 0 $X=339140 $Y=799420
X64 162 2 2036 1 INV1S $T=341000 799800 0 0 $X=341000 $Y=799420
X65 1996 2 158 1 INV1S $T=341620 850200 1 0 $X=341620 $Y=844780
X66 1892 2 2046 1 INV1S $T=342860 799800 0 0 $X=342860 $Y=799420
X67 198 2 2056 1 INV1S $T=346580 799800 0 180 $X=345340 $Y=794380
X68 1864 2 2114 1 INV1S $T=351540 789720 0 0 $X=351540 $Y=789340
X69 2073 2 151 1 INV1S $T=351540 840120 0 0 $X=351540 $Y=839740
X70 2152 2 205 1 INV1S $T=355880 759480 1 180 $X=354640 $Y=759100
X71 215 2 2157 1 INV1S $T=360220 799800 0 0 $X=360220 $Y=799420
X72 2156 2 1869 1 INV1S $T=360840 880440 0 0 $X=360840 $Y=880060
X73 2122 2 2065 1 INV1S $T=362080 860280 1 0 $X=362080 $Y=854860
X74 2151 2 1871 1 INV1S $T=363320 850200 0 0 $X=363320 $Y=849820
X75 222 2 2181 1 INV1S $T=363940 799800 0 0 $X=363940 $Y=799420
X76 2200 2 1856 1 INV1S $T=367660 870360 0 180 $X=366420 $Y=864940
X77 2206 2 153 1 INV1S $T=368280 860280 0 180 $X=367040 $Y=854860
X78 2204 2 2212 1 INV1S $T=368280 809880 1 0 $X=368280 $Y=804460
X79 1828 2 2226 1 INV1S $T=370760 830040 1 0 $X=370760 $Y=824620
X80 209 2 2236 1 INV1S $T=373860 860280 1 180 $X=372620 $Y=859900
X81 2250 2 2200 1 INV1S $T=375100 819960 1 180 $X=373860 $Y=819580
X82 226 2 1740 1 INV1S $T=375720 769560 1 180 $X=374480 $Y=769180
X83 1704 2 2257 1 INV1S $T=375100 789720 0 0 $X=375100 $Y=789340
X84 2263 2 2289 1 INV1S $T=377580 819960 1 0 $X=377580 $Y=814540
X85 217 2 252 1 INV1S $T=380060 870360 1 0 $X=380060 $Y=864940
X86 2281 2 2305 1 INV1S $T=380680 799800 1 0 $X=380680 $Y=794380
X87 2227 2 1912 1 INV1S $T=381300 850200 0 0 $X=381300 $Y=849820
X88 1886 2 172 1 INV1S $T=382540 860280 1 180 $X=381300 $Y=859900
X89 2277 2 2306 1 INV1S $T=381920 799800 0 0 $X=381920 $Y=799420
X90 2317 2 2063 1 INV1S $T=384400 840120 1 180 $X=383160 $Y=839740
X91 2177 2 255 1 INV1S $T=386260 860280 1 0 $X=386260 $Y=854860
X92 2322 2 2342 1 INV1S $T=389360 809880 0 180 $X=388120 $Y=804460
X93 2226 2 2334 1 INV1S $T=389980 830040 1 180 $X=388740 $Y=829660
X94 2370 2 1952 1 INV1S $T=391220 749400 0 180 $X=389980 $Y=743980
X95 2337 2 2360 1 INV1S $T=389980 809880 1 0 $X=389980 $Y=804460
X96 2226 2 2343 1 INV1S $T=390600 830040 0 0 $X=390600 $Y=829660
X97 2330 2 2310 1 INV1S $T=391840 870360 1 180 $X=390600 $Y=869980
X98 2303 2 2323 1 INV1S $T=393080 819960 1 0 $X=393080 $Y=814540
X99 154 2 270 1 INV1S $T=394320 890520 1 180 $X=393080 $Y=890140
X100 2367 2 2382 1 INV1S $T=394940 840120 0 180 $X=393700 $Y=834700
X101 2376 2 2385 1 INV1S $T=394320 799800 0 0 $X=394320 $Y=799420
X102 2404 2 2396 1 INV1S $T=398040 860280 0 180 $X=396800 $Y=854860
X103 2400 2 2206 1 INV1S $T=399280 819960 1 180 $X=398040 $Y=819580
X104 2161 2 2191 1 INV1S $T=399900 880440 0 0 $X=399900 $Y=880060
X105 227 2 236 1 INV1S $T=400520 880440 1 0 $X=400520 $Y=875020
X106 2399 2 2430 1 INV1S $T=403000 840120 0 0 $X=403000 $Y=839740
X107 2444 2 2447 1 INV1S $T=405480 819960 1 180 $X=404240 $Y=819580
X108 2425 2 2459 1 INV1S $T=404860 850200 0 0 $X=404860 $Y=849820
X109 292 2 2152 1 INV1S $T=409820 749400 1 180 $X=408580 $Y=749020
X110 2152 2 2465 1 INV1S $T=408580 759480 0 0 $X=408580 $Y=759100
X111 2487 2 2470 1 INV1S $T=410440 840120 1 180 $X=409200 $Y=839740
X112 2494 2 2100 1 INV1S $T=411680 850200 0 180 $X=410440 $Y=844780
X113 2476 2 235 1 INV1S $T=411060 830040 1 0 $X=411060 $Y=824620
X114 2403 2 2300 1 INV1S $T=412920 880440 0 180 $X=411680 $Y=875020
X115 2513 2 2523 1 INV1S $T=414780 819960 1 0 $X=414780 $Y=814540
X116 2554 2 2317 1 INV1S $T=423460 840120 0 180 $X=422220 $Y=834700
X117 2317 2 2571 1 INV1S $T=424080 850200 1 0 $X=424080 $Y=844780
X118 1893 2 2287 1 INV1S $T=424700 840120 1 0 $X=424700 $Y=834700
X119 2514 2 2583 1 INV1S $T=428420 860280 0 0 $X=428420 $Y=859900
X120 2420 2 269 1 INV1S $T=429660 870360 1 0 $X=429660 $Y=864940
X121 2370 2 2554 1 INV1S $T=434000 809880 1 180 $X=432760 $Y=809500
X122 2211 2 276 1 INV1S $T=435240 880440 0 0 $X=435240 $Y=880060
X123 2305 2 2630 1 INV1S $T=437100 799800 1 0 $X=437100 $Y=794380
X124 2532 2 2638 1 INV1S $T=438340 809880 0 0 $X=438340 $Y=809500
X125 2583 2 2632 1 INV1S $T=439580 860280 0 0 $X=439580 $Y=859900
X126 2638 2 2620 1 INV1S $T=442060 799800 1 180 $X=440820 $Y=799420
X127 2641 2 2649 1 INV1S $T=440820 809880 0 0 $X=440820 $Y=809500
X128 337 2 2652 1 INV1S $T=441440 870360 1 0 $X=441440 $Y=864940
X129 2655 2 2660 1 INV1S $T=443300 779640 1 0 $X=443300 $Y=774220
X130 2638 2 2697 1 INV1S $T=447020 809880 0 0 $X=447020 $Y=809500
X131 347 2 349 1 INV1S $T=450740 809880 1 0 $X=450740 $Y=804460
X132 2708 2 2712 1 INV1S $T=451360 779640 0 0 $X=451360 $Y=779260
X133 360 2 358 1 INV1S $T=458800 729240 1 180 $X=457560 $Y=728860
X134 363 2 2370 1 INV1S $T=460660 739320 1 180 $X=459420 $Y=738940
X135 2242 2 2708 1 INV1S $T=460040 769560 1 0 $X=460040 $Y=764140
X136 360 2 292 1 INV1S $T=463140 729240 1 0 $X=463140 $Y=723820
X137 2301 2 2706 1 INV1S $T=463140 779640 0 0 $X=463140 $Y=779260
X138 345 2 2785 1 INV1S $T=466240 880440 0 0 $X=466240 $Y=880060
X139 2784 2 370 1 INV1S $T=466860 870360 0 0 $X=466860 $Y=869980
X140 2801 2 2690 1 INV1S $T=469960 830040 1 180 $X=468720 $Y=829660
X141 2299 2 2784 1 INV1S $T=469960 830040 0 0 $X=469960 $Y=829660
X142 2667 2 2821 1 INV1S $T=470580 799800 1 0 $X=470580 $Y=794380
X143 2821 2 2797 1 INV1S $T=473060 809880 0 180 $X=471820 $Y=804460
X144 2785 2 2816 1 INV1S $T=473060 880440 1 180 $X=471820 $Y=880060
X145 376 2 2819 1 INV1S $T=474300 729240 0 180 $X=473060 $Y=723820
X146 2821 2 2782 1 INV1S $T=474300 799800 1 0 $X=474300 $Y=794380
X147 2833 2 363 1 INV1S $T=475540 739320 0 0 $X=475540 $Y=738940
X148 2843 2 2801 1 INV1S $T=477400 830040 1 180 $X=476160 $Y=829660
X149 387 2 377 1 INV1S $T=479880 739320 0 180 $X=478640 $Y=733900
X150 2857 2 2852 1 INV1S $T=481740 840120 1 180 $X=480500 $Y=839740
X151 2301 2 2898 1 INV1S $T=489800 749400 1 180 $X=488560 $Y=749020
X152 2849 2 402 1 INV1S $T=492900 769560 1 0 $X=492900 $Y=764140
X153 2984 2 2828 1 INV1S $T=505300 880440 1 180 $X=504060 $Y=880060
X154 2997 2 2933 1 INV1S $T=507160 769560 0 180 $X=505920 $Y=764140
X155 2952 2 399 1 INV1S $T=507780 840120 0 180 $X=506540 $Y=834700
X156 424 2 2930 1 INV1S $T=509020 809880 1 180 $X=507780 $Y=809500
X157 2580 2 2987 1 INV1S $T=508400 789720 1 0 $X=508400 $Y=784300
X158 424 2 2907 1 INV1S $T=510880 880440 1 0 $X=510880 $Y=875020
X159 2984 2 3034 1 INV1S $T=513980 870360 1 0 $X=513980 $Y=864940
X160 2907 2 2984 1 INV1S $T=513980 880440 1 0 $X=513980 $Y=875020
X161 3049 2 2947 1 INV1S $T=518940 819960 0 0 $X=518940 $Y=819580
X162 435 2 3077 1 INV1S $T=521420 840120 0 0 $X=521420 $Y=839740
X163 436 2 403 1 INV1S $T=522660 900600 0 180 $X=521420 $Y=895180
X164 3095 2 436 1 INV1S $T=527620 900600 0 180 $X=526380 $Y=895180
X165 3128 2 3060 1 INV1S $T=531340 729240 0 180 $X=530100 $Y=723820
X166 3128 2 444 1 INV1S $T=532580 729240 1 0 $X=532580 $Y=723820
X167 3168 2 2882 1 INV1S $T=536920 850200 1 180 $X=535680 $Y=849820
X168 3169 2 2999 1 INV1S $T=536920 880440 1 180 $X=535680 $Y=880060
X169 2301 2 428 1 INV1S $T=536300 749400 0 0 $X=536300 $Y=749020
X170 2306 2 3167 1 INV1S $T=536300 789720 0 0 $X=536300 $Y=789340
X171 2997 2 3149 1 INV1S $T=538780 779640 0 180 $X=537540 $Y=774220
X172 3181 2 2977 1 INV1S $T=540020 789720 0 180 $X=538780 $Y=784300
X173 2234 2 3161 1 INV1S $T=538780 789720 0 0 $X=538780 $Y=789340
X174 2785 2 3186 1 INV1S $T=538780 880440 0 0 $X=538780 $Y=880060
X175 3187 2 3093 1 INV1S $T=541880 819960 0 180 $X=540640 $Y=814540
X176 3190 2 2997 1 INV1S $T=542500 779640 0 180 $X=541260 $Y=774220
X177 3167 2 3101 1 INV1S $T=546220 830040 1 180 $X=544980 $Y=829660
X178 2306 2 3225 1 INV1S $T=549940 809880 1 0 $X=549940 $Y=804460
X179 3240 2 2965 1 INV1S $T=553660 819960 1 180 $X=552420 $Y=819580
X180 3246 2 3199 1 INV1S $T=554900 789720 1 180 $X=553660 $Y=789340
X181 3157 2 3246 1 INV1S $T=553660 799800 0 0 $X=553660 $Y=799420
X182 3246 2 3223 1 INV1S $T=554280 789720 1 0 $X=554280 $Y=784300
X183 459 2 3259 1 INV1S $T=556760 789720 1 0 $X=556760 $Y=784300
X184 3259 2 3094 1 INV1S $T=559240 819960 1 180 $X=558000 $Y=819580
X185 3259 2 3285 1 INV1S $T=561100 819960 1 0 $X=561100 $Y=814540
X186 466 2 3288 1 INV1S $T=561720 860280 1 0 $X=561720 $Y=854860
X187 3227 2 3290 1 INV1S $T=561720 860280 0 0 $X=561720 $Y=859900
X188 3288 2 3247 1 INV1S $T=562340 840120 0 0 $X=562340 $Y=839740
X189 3304 2 3298 1 INV1S $T=564820 779640 1 180 $X=563580 $Y=779260
X190 3301 2 482 1 INV1S $T=565440 809880 1 180 $X=564200 $Y=809500
X191 3304 2 3035 1 INV1S $T=564820 779640 0 0 $X=564820 $Y=779260
X192 3315 2 3304 1 INV1S $T=567300 779640 1 180 $X=566060 $Y=779260
X193 3151 2 3316 1 INV1S $T=566060 840120 1 0 $X=566060 $Y=834700
X194 3321 2 3287 1 INV1S $T=567920 860280 1 180 $X=566680 $Y=859900
X195 494 2 3328 1 INV1S $T=569160 759480 0 0 $X=569160 $Y=759100
X196 3015 2 3003 1 INV1S $T=570400 809880 0 180 $X=569160 $Y=804460
X197 3328 2 3202 1 INV1S $T=569780 759480 1 0 $X=569780 $Y=754060
X198 3263 2 3343 1 INV1S $T=572880 779640 1 180 $X=571640 $Y=779260
X199 3290 2 3397 1 INV1S $T=577220 870360 0 0 $X=577220 $Y=869980
X200 3403 2 3382 1 INV1S $T=579700 749400 1 180 $X=578460 $Y=749020
X201 3393 2 3384 1 INV1S $T=579080 799800 1 0 $X=579080 $Y=794380
X202 2234 2 3393 1 INV1S $T=579700 789720 1 0 $X=579700 $Y=784300
X203 3403 2 3413 1 INV1S $T=580940 759480 1 0 $X=580940 $Y=754060
X204 3417 2 3256 1 INV1S $T=582800 789720 0 180 $X=581560 $Y=784300
X205 3252 2 3403 1 INV1S $T=583420 749400 1 0 $X=583420 $Y=743980
X206 3420 2 3418 1 INV1S $T=584660 759480 1 180 $X=583420 $Y=759100
X207 3135 2 3420 1 INV1S $T=583420 769560 1 0 $X=583420 $Y=764140
X208 3420 2 3430 1 INV1S $T=585280 769560 1 0 $X=585280 $Y=764140
X209 2234 2 534 1 INV1S $T=588380 749400 1 0 $X=588380 $Y=743980
X210 3454 2 497 1 INV1S $T=593960 749400 0 180 $X=592720 $Y=743980
X211 3454 2 540 1 INV1S $T=593340 809880 1 0 $X=593340 $Y=804460
X212 3343 2 3407 1 INV1S $T=595820 749400 0 180 $X=594580 $Y=743980
X213 3495 2 3454 1 INV1S $T=599540 779640 1 180 $X=598300 $Y=779260
X214 529 2 545 1 INV1S $T=598920 739320 0 0 $X=598920 $Y=738940
X215 3494 2 3485 1 INV1S $T=600780 880440 0 180 $X=599540 $Y=875020
X216 3316 2 3520 1 INV1S $T=605120 840120 1 0 $X=605120 $Y=834700
X217 3352 2 3536 1 INV1S $T=609460 860280 1 180 $X=608220 $Y=859900
X218 3553 2 554 1 INV1S $T=611940 890520 0 180 $X=610700 $Y=885100
X219 3473 2 3562 1 INV1S $T=615660 809880 0 0 $X=615660 $Y=809500
X220 3428 2 3575 1 INV1S $T=615660 870360 1 0 $X=615660 $Y=864940
X221 3575 2 563 1 INV1S $T=616280 890520 1 0 $X=616280 $Y=885100
X222 3582 2 557 1 INV1S $T=617520 880440 0 0 $X=617520 $Y=880060
X223 572 2 565 1 INV1S $T=619380 729240 1 180 $X=618140 $Y=728860
X224 3575 2 3572 1 INV1S $T=618140 870360 1 0 $X=618140 $Y=864940
X225 3607 2 3490 1 INV1S $T=623100 769560 0 180 $X=621860 $Y=764140
X226 3609 2 3597 1 INV1S $T=622480 840120 1 0 $X=622480 $Y=834700
X227 3463 2 3467 1 INV1S $T=624960 769560 0 180 $X=623720 $Y=764140
X228 3487 2 3463 1 INV1S $T=623720 769560 0 0 $X=623720 $Y=769180
X229 3636 2 3510 1 INV1S $T=624960 850200 0 180 $X=623720 $Y=844780
X230 3627 2 3484 1 INV1S $T=624960 870360 1 0 $X=624960 $Y=864940
X231 3407 2 590 1 INV1S $T=627440 729240 0 0 $X=627440 $Y=728860
X232 3636 2 3592 1 INV1S $T=629300 850200 0 180 $X=628060 $Y=844780
X233 3656 2 3655 1 INV1S $T=630540 870360 0 0 $X=630540 $Y=869980
X234 577 2 3636 1 INV1S $T=633020 850200 0 180 $X=631780 $Y=844780
X235 605 2 572 1 INV1S $T=634880 729240 0 180 $X=633640 $Y=723820
X236 3673 2 3657 1 INV1S $T=635500 830040 1 180 $X=634260 $Y=829660
X237 3673 2 3555 1 INV1S $T=636740 830040 0 180 $X=635500 $Y=824620
X238 3680 2 608 1 INV1S $T=636740 880440 0 180 $X=635500 $Y=875020
X239 3552 2 3686 1 INV1S $T=636740 809880 0 0 $X=636740 $Y=809500
X240 3592 2 3673 1 INV1S $T=637980 830040 0 180 $X=636740 $Y=824620
X241 2301 2 3692 1 INV1S $T=637980 769560 0 0 $X=637980 $Y=769180
X242 618 2 615 1 INV1S $T=640460 729240 0 180 $X=639220 $Y=723820
X243 618 2 3544 1 INV1S $T=640460 729240 1 0 $X=640460 $Y=723820
X244 3707 2 3679 1 INV1S $T=642940 799800 1 0 $X=642940 $Y=794380
X245 3724 2 3737 1 INV1S $T=646040 850200 1 0 $X=646040 $Y=844780
X246 3729 2 3724 1 INV1S $T=647280 870360 0 180 $X=646040 $Y=864940
X247 3734 2 3519 1 INV1S $T=647900 739320 1 180 $X=646660 $Y=738940
X248 3734 2 3641 1 INV1S $T=648520 739320 0 0 $X=648520 $Y=738940
X249 3755 2 3637 1 INV1S $T=652860 799800 0 180 $X=651620 $Y=794380
X250 3761 2 3755 1 INV1S $T=653480 799800 1 0 $X=653480 $Y=794380
X251 3771 2 3687 1 INV1S $T=654720 880440 0 180 $X=653480 $Y=875020
X252 3779 2 3734 1 INV1S $T=657200 739320 1 180 $X=655960 $Y=738940
X253 645 2 3667 1 INV1S $T=655960 890520 0 0 $X=655960 $Y=890140
X254 3771 2 3742 1 INV1S $T=656580 860280 1 0 $X=656580 $Y=854860
X255 3755 2 3785 1 INV1S $T=657200 799800 1 0 $X=657200 $Y=794380
X256 3667 2 3771 1 INV1S $T=659680 880440 1 180 $X=658440 $Y=880060
X257 2849 2 3794 1 INV1S $T=659060 749400 1 0 $X=659060 $Y=743980
X258 3803 2 3729 1 INV1S $T=660920 870360 1 180 $X=659680 $Y=869980
X259 3773 2 656 1 INV1S $T=662160 880440 1 0 $X=662160 $Y=875020
X260 659 2 577 1 INV1S $T=665260 830040 0 180 $X=664020 $Y=824620
X261 3697 2 663 1 INV1S $T=668360 890520 1 180 $X=667120 $Y=890140
X262 3836 2 3825 1 INV1S $T=669600 880440 0 180 $X=668360 $Y=875020
X263 3892 2 3800 1 INV1S $T=678900 789720 0 180 $X=677660 $Y=784300
X264 3892 2 3881 1 INV1S $T=679520 779640 0 0 $X=679520 $Y=779260
X265 3887 2 3892 1 INV1S $T=681380 799800 0 180 $X=680140 $Y=794380
X266 3900 2 3858 1 INV1S $T=681380 870360 0 180 $X=680140 $Y=864940
X267 659 2 3887 1 INV1S $T=682000 819960 0 180 $X=680760 $Y=814540
X268 3903 2 698 1 INV1S $T=685720 890520 0 0 $X=685720 $Y=890140
X269 3956 2 3900 1 INV1S $T=691300 870360 0 180 $X=690060 $Y=864940
X270 3972 2 692 1 INV1S $T=693160 880440 0 180 $X=691920 $Y=875020
X271 3981 2 3864 1 INV1S $T=695640 729240 1 180 $X=694400 $Y=728860
X272 719 2 3981 1 INV1S $T=698740 729240 1 180 $X=697500 $Y=728860
X273 3981 2 3779 1 INV1S $T=697500 739320 1 0 $X=697500 $Y=733900
X274 3859 2 4057 1 INV1S $T=706180 860280 1 0 $X=706180 $Y=854860
X275 4034 2 4029 1 INV1S $T=706800 779640 1 0 $X=706800 $Y=774220
X276 4101 2 4050 1 INV1S $T=713620 870360 1 180 $X=712380 $Y=869980
X277 4104 2 3947 1 INV1S $T=714860 779640 0 180 $X=713620 $Y=774220
X278 4112 2 685 1 INV1S $T=715480 729240 1 180 $X=714240 $Y=728860
X279 4146 2 3828 1 INV1S $T=722300 789720 1 180 $X=721060 $Y=789340
X280 4144 2 4136 1 INV1S $T=721060 830040 0 0 $X=721060 $Y=829660
X281 4148 2 757 1 INV1S $T=722920 729240 0 180 $X=721680 $Y=723820
X282 4155 2 3906 1 INV1S $T=724160 749400 1 180 $X=722920 $Y=749020
X283 3211 2 4161 1 INV1S $T=722920 789720 0 0 $X=722920 $Y=789340
X284 4170 2 3867 1 INV1S $T=728500 769560 1 180 $X=727260 $Y=769180
X285 4173 2 3822 1 INV1S $T=729120 739320 0 180 $X=727880 $Y=733900
X286 4161 2 4130 1 INV1S $T=729120 789720 1 180 $X=727880 $Y=789340
X287 4057 2 4167 1 INV1S $T=730360 860280 0 180 $X=729120 $Y=854860
X288 4161 2 3994 1 INV1S $T=730980 809880 1 180 $X=729740 $Y=809500
X289 777 2 4185 1 INV1S $T=730980 789720 1 0 $X=730980 $Y=784300
X290 4012 2 4179 1 INV1S $T=730980 789720 0 0 $X=730980 $Y=789340
X291 4204 2 4127 1 INV1S $T=732840 840120 1 180 $X=731600 $Y=839740
X292 774 2 4181 1 INV1S $T=734080 759480 0 180 $X=732840 $Y=754060
X293 4191 2 4183 1 INV1S $T=734080 769560 0 180 $X=732840 $Y=764140
X294 4195 2 460 1 INV1S $T=734080 779640 1 180 $X=732840 $Y=779260
X295 4161 2 4178 1 INV1S $T=734700 819960 1 0 $X=734700 $Y=814540
X296 788 2 787 1 INV1S $T=736560 799800 0 180 $X=735320 $Y=794380
X297 4218 2 765 1 INV1S $T=737800 779640 1 180 $X=736560 $Y=779260
X298 4219 2 789 1 INV1S $T=737800 799800 0 180 $X=736560 $Y=794380
X299 4225 2 3507 1 INV1S $T=738420 769560 1 180 $X=737180 $Y=769180
X300 4242 2 4208 1 INV1S $T=740900 739320 0 180 $X=739660 $Y=733900
X301 4241 2 772 1 INV1S $T=740900 789720 1 180 $X=739660 $Y=789340
X302 4236 2 4176 1 INV1S $T=739660 819960 1 0 $X=739660 $Y=814540
X303 659 2 4224 1 INV1S $T=740280 799800 1 0 $X=740280 $Y=794380
X304 805 2 4162 1 INV1S $T=742140 749400 0 180 $X=740900 $Y=743980
X305 4246 2 803 1 INV1S $T=742760 789720 1 180 $X=741520 $Y=789340
X306 4267 2 813 1 INV1S $T=745860 789720 0 0 $X=745860 $Y=789340
X307 4272 2 819 1 INV1S $T=747720 779640 0 0 $X=747720 $Y=779260
X308 4282 2 458 1 INV1S $T=748960 789720 1 180 $X=747720 $Y=789340
X309 4290 2 823 1 INV1S $T=751440 799800 1 180 $X=750200 $Y=799420
X310 4294 2 825 1 INV1S $T=752060 789720 0 180 $X=750820 $Y=784300
X311 4288 2 776 1 INV1S $T=751440 779640 1 0 $X=751440 $Y=774220
X312 4289 2 826 1 INV1S $T=751440 789720 0 0 $X=751440 $Y=789340
X313 4303 2 788 1 INV1S $T=753920 779640 1 180 $X=752680 $Y=779260
X314 4310 2 827 1 INV1S $T=755160 789720 0 180 $X=753920 $Y=784300
X315 4309 2 3532 1 INV1S $T=755780 739320 1 0 $X=755780 $Y=733900
X316 4322 2 4234 1 INV1S $T=756400 840120 1 0 $X=756400 $Y=834700
X317 4327 2 805 1 INV1S $T=758880 769560 1 180 $X=757640 $Y=769180
X318 4178 2 833 1 INV1S $T=757640 850200 0 0 $X=757640 $Y=849820
X319 832 2 4302 1 INV1S $T=758880 729240 1 0 $X=758880 $Y=723820
X320 4276 2 4300 1 INV1S $T=758880 769560 0 0 $X=758880 $Y=769180
X321 4348 2 799 1 INV1S $T=762600 769560 0 180 $X=761360 $Y=764140
X322 4326 2 4347 1 INV1S $T=765700 729240 0 0 $X=765700 $Y=728860
X323 4383 2 4359 1 INV1S $T=768180 890520 1 180 $X=766940 $Y=890140
X324 4266 2 4385 1 INV1S $T=767560 850200 1 0 $X=767560 $Y=844780
X325 4374 2 4383 1 INV1S $T=768180 890520 1 0 $X=768180 $Y=885100
X326 4387 2 4384 1 INV1S $T=769420 749400 0 0 $X=769420 $Y=749020
X327 4388 2 4380 1 INV1S $T=770040 769560 1 0 $X=770040 $Y=764140
X328 4393 2 4360 1 INV1S $T=771280 809880 1 180 $X=770040 $Y=809500
X329 4409 2 4400 1 INV1S $T=773760 809880 1 180 $X=772520 $Y=809500
X330 4409 2 861 1 INV1S $T=774380 850200 1 180 $X=773140 $Y=849820
X331 4424 2 4374 1 INV1S $T=774380 860280 0 180 $X=773140 $Y=854860
X332 4439 2 4352 1 INV1S $T=776860 890520 0 180 $X=775620 $Y=885100
X333 4450 2 4393 1 INV1S $T=778720 819960 0 180 $X=777480 $Y=814540
X334 4378 2 4463 1 INV1S $T=779960 729240 0 0 $X=779960 $Y=728860
X335 4349 2 4517 1 INV1S $T=791740 789720 1 180 $X=790500 $Y=789340
X336 4555 2 4512 1 INV1S $T=796700 850200 1 180 $X=795460 $Y=849820
X337 4564 2 4491 1 INV1S $T=797320 870360 0 180 $X=796080 $Y=864940
X338 4495 2 4499 1 INV1S $T=799800 840120 1 0 $X=799800 $Y=834700
X339 4581 2 4578 1 INV1S $T=801660 779640 1 180 $X=800420 $Y=779260
X340 4454 2 906 1 INV1S $T=800420 890520 0 0 $X=800420 $Y=890140
X341 4495 2 4589 1 INV1S $T=801040 799800 1 0 $X=801040 $Y=794380
X342 4454 2 4590 1 INV1S $T=801040 880440 1 0 $X=801040 $Y=875020
X343 4596 2 4600 1 INV1S $T=802280 870360 0 0 $X=802280 $Y=869980
X344 4605 2 4596 1 INV1S $T=804760 870360 1 180 $X=803520 $Y=869980
X345 4434 2 928 1 INV1S $T=805380 729240 0 0 $X=805380 $Y=728860
X346 888 2 4361 1 INV1S $T=806620 830040 1 180 $X=805380 $Y=829660
X347 4600 2 4544 1 INV1S $T=805380 890520 0 0 $X=805380 $Y=890140
X348 925 2 924 1 INV1S $T=807860 729240 0 180 $X=806620 $Y=723820
X349 4578 2 4628 1 INV1S $T=807240 789720 0 0 $X=807240 $Y=789340
X350 4600 2 887 1 INV1S $T=808480 890520 1 0 $X=808480 $Y=885100
X351 4642 2 4608 1 INV1S $T=810340 779640 1 180 $X=809100 $Y=779260
X352 4643 2 4648 1 INV1S $T=809720 789720 0 0 $X=809720 $Y=789340
X353 4589 2 4650 1 INV1S $T=810960 799800 1 0 $X=810960 $Y=794380
X354 4656 2 4585 1 INV1S $T=812820 759480 1 0 $X=812820 $Y=754060
X355 4431 2 4662 1 INV1S $T=813440 749400 1 0 $X=813440 $Y=743980
X356 4266 2 931 1 INV1S $T=815920 880440 0 180 $X=814680 $Y=875020
X357 4683 2 4505 1 INV1S $T=817780 809880 1 180 $X=816540 $Y=809500
X358 4704 2 4645 1 INV1S $T=820880 729240 1 0 $X=820880 $Y=723820
X359 4706 2 4716 1 INV1S $T=820880 870360 0 0 $X=820880 $Y=869980
X360 4707 2 941 1 INV1S $T=820880 890520 0 0 $X=820880 $Y=890140
X361 4734 2 4728 1 INV1S $T=826460 759480 0 180 $X=825220 $Y=754060
X362 4639 2 4734 1 INV1S $T=825840 769560 1 0 $X=825840 $Y=764140
X363 848 2 4707 1 INV1S $T=826460 880440 0 0 $X=826460 $Y=880060
X364 4736 2 948 1 INV1S $T=827700 900600 0 180 $X=826460 $Y=895180
X365 4755 2 951 1 INV1S $T=829560 850200 1 180 $X=828320 $Y=849820
X366 4721 2 4755 1 INV1S $T=830800 840120 1 0 $X=830800 $Y=834700
X367 4777 2 4683 1 INV1S $T=833280 799800 0 180 $X=832040 $Y=794380
X368 4487 2 4780 1 INV1S $T=832660 789720 0 0 $X=832660 $Y=789340
X369 4789 2 4699 1 INV1S $T=835140 749400 0 180 $X=833900 $Y=743980
X370 4683 2 4785 1 INV1S $T=833900 799800 1 0 $X=833900 $Y=794380
X371 4755 2 4791 1 INV1S $T=835760 840120 0 0 $X=835760 $Y=839740
X372 4734 2 4806 1 INV1S $T=837000 749400 0 0 $X=837000 $Y=749020
X373 4734 2 4725 1 INV1S $T=837620 759480 0 0 $X=837620 $Y=759100
X374 4813 2 4712 1 INV1S $T=838860 850200 1 180 $X=837620 $Y=849820
X375 4707 2 4815 1 INV1S $T=839480 900600 1 0 $X=839480 $Y=895180
X376 4810 2 4821 1 INV1S $T=840100 799800 1 0 $X=840100 $Y=794380
X377 4833 2 4824 1 INV1S $T=843820 830040 1 180 $X=842580 $Y=829660
X378 4839 2 4813 1 INV1S $T=845060 850200 0 180 $X=843820 $Y=844780
X379 4813 2 4852 1 INV1S $T=845060 850200 1 0 $X=845060 $Y=844780
X380 4795 2 4866 1 INV1S $T=846300 779640 0 0 $X=846300 $Y=779260
X381 973 2 4839 1 INV1S $T=848780 850200 0 180 $X=847540 $Y=844780
X382 4780 2 4871 1 INV1S $T=848160 789720 0 0 $X=848160 $Y=789340
X383 4876 2 4814 1 INV1S $T=851880 840120 0 180 $X=850640 $Y=834700
X384 4878 2 4439 1 INV1S $T=851260 880440 0 0 $X=851260 $Y=880060
X385 4666 2 4902 1 INV1S $T=853740 819960 1 0 $X=853740 $Y=814540
X386 4700 2 4833 1 INV1S $T=853740 830040 1 0 $X=853740 $Y=824620
X387 4895 2 4731 1 INV1S $T=854360 860280 1 0 $X=854360 $Y=854860
X388 4815 2 4901 1 INV1S $T=854360 900600 1 0 $X=854360 $Y=895180
X389 973 2 980 1 INV1S $T=858700 890520 1 0 $X=858700 $Y=885100
X390 4383 2 985 1 INV1S $T=865520 890520 1 0 $X=865520 $Y=885100
X391 4902 2 1003 1 INV1S $T=879780 890520 1 0 $X=879780 $Y=885100
X392 4902 2 5030 1 INV1S $T=880400 819960 1 0 $X=880400 $Y=814540
X393 5100 2 4975 1 INV1S $T=892180 809880 1 180 $X=890940 $Y=809500
X394 5100 2 5096 1 INV1S $T=892180 819960 0 180 $X=890940 $Y=814540
X395 1026 2 5100 1 INV1S $T=897760 819960 0 180 $X=896520 $Y=814540
X396 4439 2 1030 1 INV1S $T=899620 890520 0 0 $X=899620 $Y=890140
X397 4353 2 5162 1 INV1S $T=902100 769560 1 0 $X=902100 $Y=764140
X398 990 2 5178 1 INV1S $T=903340 900600 1 0 $X=903340 $Y=895180
X399 5177 2 5212 1 INV1S $T=908920 769560 0 0 $X=908920 $Y=769180
X400 5178 2 5191 1 INV1S $T=910780 900600 1 0 $X=910780 $Y=895180
X401 5248 2 5181 1 INV1S $T=918840 809880 0 180 $X=917600 $Y=804460
X402 5178 2 1044 1 INV1S $T=917600 900600 1 0 $X=917600 $Y=895180
X403 5231 2 5233 1 INV1S $T=918220 779640 0 0 $X=918220 $Y=779260
X404 5248 2 5253 1 INV1S $T=921320 809880 1 0 $X=921320 $Y=804460
X405 5242 2 5248 1 INV1S $T=922560 809880 1 180 $X=921320 $Y=809500
X406 5244 2 5256 1 INV1S $T=921940 840120 0 0 $X=921940 $Y=839740
X407 5250 2 5260 1 INV1S $T=923180 799800 1 0 $X=923180 $Y=794380
X408 5252 2 5267 1 INV1S $T=925040 769560 0 0 $X=925040 $Y=769180
X409 5262 2 5269 1 INV1S $T=925660 860280 1 0 $X=925660 $Y=854860
X410 5288 2 5285 1 INV1S $T=929380 870360 0 180 $X=928140 $Y=864940
X411 5288 2 5297 1 INV1S $T=933100 870360 1 180 $X=931860 $Y=869980
X412 5325 2 5288 1 INV1S $T=934340 870360 1 180 $X=933100 $Y=869980
X413 5331 2 5325 1 INV1S $T=935580 870360 1 180 $X=934340 $Y=869980
X414 5319 2 1056 1 INV1S $T=936200 830040 0 0 $X=936200 $Y=829660
X415 1058 2 5354 1 INV1S $T=938060 880440 1 0 $X=938060 $Y=875020
X416 5260 2 5374 1 INV1S $T=940540 789720 0 0 $X=940540 $Y=789340
X417 5374 2 5280 1 INV1S $T=943020 769560 0 180 $X=941780 $Y=764140
X418 5374 2 5379 1 INV1S $T=942400 789720 0 0 $X=942400 $Y=789340
X419 5380 2 5316 1 INV1S $T=943020 799800 1 0 $X=943020 $Y=794380
X420 5391 2 5286 1 INV1S $T=944880 739320 1 180 $X=943640 $Y=738940
X421 5267 2 5391 1 INV1S $T=944260 779640 1 0 $X=944260 $Y=774220
X422 5391 2 5393 1 INV1S $T=944880 739320 0 0 $X=944880 $Y=738940
X423 5309 2 5380 1 INV1S $T=944880 759480 0 0 $X=944880 $Y=759100
X424 5411 2 5293 1 INV1S $T=947980 850200 0 180 $X=946740 $Y=844780
X425 5380 2 5356 1 INV1S $T=947980 799800 1 0 $X=947980 $Y=794380
X426 5356 2 5411 1 INV1S $T=950460 850200 1 0 $X=950460 $Y=844780
X427 5385 2 5494 1 INV1S $T=960380 789720 1 0 $X=960380 $Y=784300
X428 5494 2 5307 1 INV1S $T=961620 819960 1 0 $X=961620 $Y=814540
X429 5431 2 1067 1 INV1S $T=963480 850200 1 0 $X=963480 $Y=844780
X430 5590 2 5384 1 INV1S $T=976500 850200 0 180 $X=975260 $Y=844780
X431 1103 2 1104 1 INV1S $T=980220 729240 1 0 $X=980220 $Y=723820
X432 5640 2 5590 1 INV1S $T=988280 850200 1 180 $X=987040 $Y=849820
X433 1107 2 5638 1 INV1S $T=988280 870360 1 180 $X=987040 $Y=869980
X434 5638 2 5640 1 INV1S $T=987040 880440 1 0 $X=987040 $Y=875020
X435 5590 2 5651 1 INV1S $T=990140 850200 0 0 $X=990140 $Y=849820
X436 5667 2 1110 1 INV1S $T=993240 779640 0 180 $X=992000 $Y=774220
X437 5590 2 5657 1 INV1S $T=992000 850200 0 0 $X=992000 $Y=849820
X438 5655 2 5659 1 INV1S $T=992000 860280 0 0 $X=992000 $Y=859900
X439 1114 2 5667 1 INV1S $T=998200 749400 0 180 $X=996960 $Y=743980
X440 5697 2 5686 1 INV1S $T=1000060 840120 1 180 $X=998820 $Y=839740
X441 5703 2 1119 1 INV1S $T=1000680 860280 1 0 $X=1000680 $Y=854860
X442 5711 2 5720 1 INV1S $T=1001920 769560 1 0 $X=1001920 $Y=764140
X443 5649 2 5703 1 INV1S $T=1002540 860280 1 0 $X=1002540 $Y=854860
X444 5729 2 5733 1 INV1S $T=1003780 789720 0 0 $X=1003780 $Y=789340
X445 5746 2 5714 1 INV1S $T=1006260 880440 0 180 $X=1005020 $Y=875020
X446 5659 2 5764 1 INV1S $T=1007500 850200 0 0 $X=1007500 $Y=849820
X447 5764 2 5781 1 INV1S $T=1009980 850200 1 0 $X=1009980 $Y=844780
X448 5782 2 5697 1 INV1S $T=1011840 840120 0 180 $X=1010600 $Y=834700
X449 1140 2 5698 1 INV1S $T=1011840 890520 1 180 $X=1010600 $Y=890140
X450 5746 2 5724 1 INV1S $T=1013700 880440 1 180 $X=1012460 $Y=880060
X451 5764 2 5797 1 INV1S $T=1013700 830040 1 0 $X=1013700 $Y=824620
X452 5794 2 5746 1 INV1S $T=1014940 880440 0 180 $X=1013700 $Y=875020
X453 5671 2 5800 1 INV1S $T=1014940 809880 0 0 $X=1014940 $Y=809500
X454 5782 2 5802 1 INV1S $T=1015560 840120 1 0 $X=1015560 $Y=834700
X455 5689 2 5829 1 INV1S $T=1021140 880440 0 0 $X=1021140 $Y=880060
X456 5703 2 5845 1 INV1S $T=1023620 860280 1 0 $X=1023620 $Y=854860
X457 5829 2 5840 1 INV1S $T=1024240 880440 0 0 $X=1024240 $Y=880060
X458 5849 2 1145 1 INV1S $T=1024860 890520 0 0 $X=1024860 $Y=890140
X459 1118 2 5868 1 INV1S $T=1026100 729240 1 0 $X=1026100 $Y=723820
X460 5800 2 5826 1 INV1S $T=1027340 809880 1 180 $X=1026100 $Y=809500
X461 5868 2 5830 1 INV1S $T=1027960 729240 1 0 $X=1027960 $Y=723820
X462 5874 2 5856 1 INV1S $T=1029820 809880 1 180 $X=1028580 $Y=809500
X463 5802 2 5875 1 INV1S $T=1028580 850200 0 0 $X=1028580 $Y=849820
X464 5869 2 5666 1 INV1S $T=1028580 880440 0 0 $X=1028580 $Y=880060
X465 5874 2 5805 1 INV1S $T=1030440 799800 1 180 $X=1029200 $Y=799420
X466 5665 2 5881 1 INV1S $T=1029820 789720 0 0 $X=1029820 $Y=789340
X467 5881 2 5870 1 INV1S $T=1032920 799800 0 180 $X=1031680 $Y=794380
X468 5891 2 5902 1 INV1S $T=1032920 860280 1 0 $X=1032920 $Y=854860
X469 5904 2 1140 1 INV1S $T=1032920 890520 0 0 $X=1032920 $Y=890140
X470 1152 2 5873 1 INV1S $T=1036020 880440 1 180 $X=1034780 $Y=880060
X471 5681 2 1176 1 INV1S $T=1038500 769560 1 0 $X=1038500 $Y=764140
X472 5800 2 5955 1 INV1S $T=1039740 809880 0 0 $X=1039740 $Y=809500
X473 5716 2 5964 1 INV1S $T=1042840 739320 0 0 $X=1042840 $Y=738940
X474 5675 2 1184 1 INV1S $T=1042840 850200 0 0 $X=1042840 $Y=849820
X475 5935 2 5972 1 INV1S $T=1044080 749400 0 0 $X=1044080 $Y=749020
X476 5972 2 5939 1 INV1S $T=1045320 759480 1 0 $X=1045320 $Y=754060
X477 5943 2 5874 1 INV1S $T=1048420 809880 1 180 $X=1047180 $Y=809500
X478 5964 2 5946 1 INV1S $T=1048420 739320 1 0 $X=1048420 $Y=733900
X479 5839 2 6023 1 INV1S $T=1054000 809880 0 0 $X=1054000 $Y=809500
X480 5964 2 6072 1 INV1S $T=1061440 729240 0 0 $X=1061440 $Y=728860
X481 1145 2 6110 1 INV1S $T=1070120 900600 1 0 $X=1070120 $Y=895180
X482 6116 2 6033 1 INV1S $T=1071980 809880 1 180 $X=1070740 $Y=809500
X483 6023 2 6108 1 INV1S $T=1070740 819960 1 0 $X=1070740 $Y=814540
X484 6003 2 6116 1 INV1S $T=1070740 819960 0 0 $X=1070740 $Y=819580
X485 6110 2 1201 1 INV1S $T=1072600 900600 0 180 $X=1071360 $Y=895180
X486 1176 2 5998 1 INV1S $T=1072600 880440 1 0 $X=1072600 $Y=875020
X487 6116 2 6123 1 INV1S $T=1073220 809880 0 0 $X=1073220 $Y=809500
X488 6110 2 1205 1 INV1S $T=1073220 900600 1 0 $X=1073220 $Y=895180
X489 5924 2 6168 1 INV1S $T=1082520 759480 0 0 $X=1082520 $Y=759100
X490 6162 2 6218 1 INV1S $T=1091820 880440 1 0 $X=1091820 $Y=875020
X491 6098 2 6253 1 INV1S $T=1097400 819960 1 0 $X=1097400 $Y=814540
X492 6253 2 6226 1 INV1S $T=1100500 830040 1 0 $X=1100500 $Y=824620
X493 6218 2 1236 1 INV1S $T=1100500 880440 0 0 $X=1100500 $Y=880060
X494 1256 2 1257 1 INV1S $T=1128400 880440 0 0 $X=1128400 $Y=880060
X495 3 1 2 6 BUF1S $T=220720 830040 0 0 $X=220720 $Y=829660
X496 20 1 2 1373 BUF1S $T=233740 759480 1 180 $X=231260 $Y=759100
X497 1408 1 2 1384 BUF1S $T=234360 779640 0 180 $X=231880 $Y=774220
X498 36 1 2 1407 BUF1S $T=237460 749400 1 180 $X=234980 $Y=749020
X499 1421 1 2 1411 BUF1S $T=236220 779640 1 0 $X=236220 $Y=774220
X500 29 1 2 1390 BUF1S $T=241180 779640 1 180 $X=238700 $Y=779260
X501 1429 1 2 42 BUF1S $T=245520 880440 1 0 $X=245520 $Y=875020
X502 1429 1 2 1512 BUF1S $T=250480 860280 0 0 $X=250480 $Y=859900
X503 50 1 2 1400 BUF1S $T=254820 759480 1 180 $X=252340 $Y=759100
X504 44 1 2 1493 BUF1S $T=257920 749400 0 0 $X=257920 $Y=749020
X505 59 1 2 62 BUF1S $T=259780 830040 1 0 $X=259780 $Y=824620
X506 1520 1 2 80 BUF1S $T=260400 840120 0 0 $X=260400 $Y=839740
X507 1580 1 2 45 BUF1S $T=264120 860280 1 180 $X=261640 $Y=859900
X508 1562 1 2 41 BUF1S $T=264740 890520 1 180 $X=262260 $Y=890140
X509 1608 1 2 1487 BUF1S $T=267840 850200 0 180 $X=265360 $Y=844780
X510 1610 1 2 1537 BUF1S $T=269080 830040 0 180 $X=266600 $Y=824620
X511 1599 1 2 1483 BUF1S $T=270940 860280 0 180 $X=268460 $Y=854860
X512 1453 1 2 74 BUF1S $T=268460 890520 0 0 $X=268460 $Y=890140
X513 1638 1 2 1409 BUF1S $T=272800 789720 1 180 $X=270320 $Y=789340
X514 1615 1 2 1548 BUF1S $T=272800 830040 0 180 $X=270320 $Y=824620
X515 75 1 2 1371 BUF1S $T=274660 729240 1 180 $X=272180 $Y=728860
X516 85 1 2 1655 BUF1S $T=279000 729240 1 0 $X=279000 $Y=723820
X517 1678 1 2 86 BUF1S $T=282100 860280 0 180 $X=279620 $Y=854860
X518 88 1 2 1644 BUF1S $T=280860 739320 1 0 $X=280860 $Y=733900
X519 92 1 2 89 BUF1S $T=283960 799800 1 180 $X=281480 $Y=799420
X520 1652 1 2 100 BUF1S $T=287680 860280 0 0 $X=287680 $Y=859900
X521 1685 1 2 101 BUF1S $T=287680 890520 1 0 $X=287680 $Y=885100
X522 1714 1 2 1608 BUF1S $T=292640 830040 1 180 $X=290160 $Y=829660
X523 1738 1 2 95 BUF1S $T=292640 890520 1 180 $X=290160 $Y=890140
X524 1752 1 2 104 BUF1S $T=294500 880440 1 180 $X=292020 $Y=880060
X525 35 1 2 1562 BUF1S $T=294500 870360 1 0 $X=294500 $Y=864940
X526 1714 1 2 1824 BUF1S $T=300700 819960 0 0 $X=300700 $Y=819580
X527 1828 1 2 1610 BUF1S $T=307520 830040 0 180 $X=305040 $Y=824620
X528 1829 1 2 1708 BUF1S $T=307520 840120 0 180 $X=305040 $Y=834700
X529 1824 1 2 75 BUF1S $T=307520 759480 1 0 $X=307520 $Y=754060
X530 1843 1 2 1615 BUF1S $T=310000 830040 0 180 $X=307520 $Y=824620
X531 1844 1 2 1721 BUF1S $T=310000 840120 0 180 $X=307520 $Y=834700
X532 1857 1 2 121 BUF1S $T=311860 890520 0 180 $X=309380 $Y=885100
X533 1796 1 2 128 BUF1S $T=313720 900600 1 0 $X=313720 $Y=895180
X534 1886 1 2 145 BUF1S $T=318680 880440 1 180 $X=316200 $Y=880060
X535 151 1 2 146 BUF1S $T=319920 900600 0 180 $X=317440 $Y=895180
X536 158 1 2 117 BUF1S $T=323640 900600 0 180 $X=321160 $Y=895180
X537 1912 1 2 1857 BUF1S $T=324880 880440 1 180 $X=322400 $Y=880060
X538 1911 1 2 122 BUF1S $T=326120 890520 0 180 $X=323640 $Y=885100
X539 1849 1 2 161 BUF1S $T=323640 900600 1 0 $X=323640 $Y=895180
X540 1921 1 2 111 BUF1S $T=325500 890520 0 0 $X=325500 $Y=890140
X541 1921 1 2 1908 BUF1S $T=327980 890520 1 0 $X=327980 $Y=885100
X542 1512 1 2 175 BUF1S $T=330460 890520 1 0 $X=330460 $Y=885100
X543 1970 1 2 1873 BUF1S $T=333560 830040 1 180 $X=331080 $Y=829660
X544 1829 1 2 1945 BUF1S $T=334180 819960 0 0 $X=334180 $Y=819580
X545 1996 1 2 127 BUF1S $T=336660 850200 0 180 $X=334180 $Y=844780
X546 1844 1 2 1942 BUF1S $T=334800 840120 0 0 $X=334800 $Y=839740
X547 116 1 2 188 BUF1S $T=336040 900600 1 0 $X=336040 $Y=895180
X548 190 1 2 1828 BUF1S $T=340380 830040 1 180 $X=337900 $Y=829660
X549 2063 1 2 1844 BUF1S $T=344100 840120 1 180 $X=341620 $Y=839740
X550 1843 1 2 2058 BUF1S $T=342240 830040 0 0 $X=342240 $Y=829660
X551 1970 1 2 2054 BUF1S $T=346580 830040 1 0 $X=346580 $Y=824620
X552 205 1 2 2084 BUF1S $T=352780 759480 1 180 $X=350300 $Y=759100
X553 1856 1 2 2156 BUF1S $T=358980 870360 1 0 $X=358980 $Y=864940
X554 213 1 2 2168 BUF1S $T=360840 729240 0 0 $X=360840 $Y=728860
X555 1855 1 2 2177 BUF1S $T=362080 860280 0 0 $X=362080 $Y=859900
X556 231 1 2 2184 BUF1S $T=368900 729240 1 180 $X=366420 $Y=728860
X557 235 1 2 129 BUF1S $T=370760 890520 0 180 $X=368280 $Y=885100
X558 2209 1 2 2113 BUF1S $T=372000 779640 0 180 $X=369520 $Y=774220
X559 2054 1 2 2164 BUF1S $T=370140 819960 0 0 $X=370140 $Y=819580
X560 2054 1 2 2182 BUF1S $T=370140 830040 0 0 $X=370140 $Y=829660
X561 2236 1 2 238 BUF1S $T=374480 890520 0 180 $X=372000 $Y=885100
X562 2227 1 2 243 BUF1S $T=376960 860280 1 180 $X=374480 $Y=859900
X563 250 1 2 2255 BUF1S $T=379440 729240 0 180 $X=376960 $Y=723820
X564 254 1 2 2121 BUF1S $T=384400 739320 0 180 $X=381920 $Y=733900
X565 1886 1 2 2311 BUF1S $T=381920 870360 1 0 $X=381920 $Y=864940
X566 2330 1 2 149 BUF1S $T=386260 890520 0 180 $X=383780 $Y=885100
X567 2310 1 2 114 BUF1S $T=389980 890520 1 180 $X=387500 $Y=890140
X568 2058 1 2 2325 BUF1S $T=390600 830040 1 0 $X=390600 $Y=824620
X569 2182 1 2 2373 BUF1S $T=390600 860280 1 0 $X=390600 $Y=854860
X570 275 1 2 2150 BUF1S $T=397420 739320 0 180 $X=394940 $Y=733900
X571 2397 1 2 154 BUF1S $T=397420 880440 1 180 $X=394940 $Y=880060
X572 2413 1 2 213 BUF1S $T=400520 739320 0 180 $X=398040 $Y=733900
X573 1912 1 2 280 BUF1S $T=398040 890520 0 0 $X=398040 $Y=890140
X574 279 1 2 2125 BUF1S $T=399900 729240 0 0 $X=399900 $Y=728860
X575 287 1 2 261 BUF1S $T=407960 729240 1 180 $X=405480 $Y=728860
X576 291 1 2 2438 BUF1S $T=410440 729240 1 180 $X=407960 $Y=728860
X577 2468 1 2 2209 BUF1S $T=412300 779640 1 0 $X=412300 $Y=774220
X578 2373 1 2 2514 BUF1S $T=412300 860280 1 0 $X=412300 $Y=854860
X579 297 1 2 2489 BUF1S $T=412920 729240 1 0 $X=412920 $Y=723820
X580 298 1 2 2468 BUF1S $T=416640 759480 0 180 $X=414160 $Y=754060
X581 2506 1 2 1796 BUF1S $T=416640 860280 1 180 $X=414160 $Y=859900
X582 2191 1 2 290 BUF1S $T=416640 890520 1 180 $X=414160 $Y=890140
X583 2546 1 2 2007 BUF1S $T=418500 840120 0 180 $X=416020 $Y=834700
X584 301 1 2 2451 BUF1S $T=419740 759480 0 180 $X=417260 $Y=754060
X585 2413 1 2 2456 BUF1S $T=424080 759480 0 180 $X=421600 $Y=754060
X586 2546 1 2 2522 BUF1S $T=424700 860280 1 180 $X=422220 $Y=859900
X587 1940 1 2 2546 BUF1S $T=425940 840120 1 0 $X=425940 $Y=834700
X588 2571 1 2 2530 BUF1S $T=429660 870360 0 180 $X=427180 $Y=864940
X589 2171 1 2 259 BUF1S $T=429660 880440 1 180 $X=427180 $Y=880060
X590 2164 1 2 2532 BUF1S $T=428420 819960 0 0 $X=428420 $Y=819580
X591 320 1 2 2474 BUF1S $T=432140 729240 0 180 $X=429660 $Y=723820
X592 353 1 2 2413 BUF1S $T=453840 739320 0 180 $X=451360 $Y=733900
X593 2708 1 2 347 BUF1S $T=451980 809880 1 0 $X=451980 $Y=804460
X594 2684 1 2 368 BUF1S $T=463760 870360 1 0 $X=463760 $Y=864940
X595 371 1 2 356 BUF1S $T=468100 890520 0 180 $X=465620 $Y=885100
X596 2828 1 2 2710 BUF1S $T=474920 870360 1 180 $X=472440 $Y=869980
X597 2828 1 2 2725 BUF1S $T=477400 850200 1 180 $X=474920 $Y=849820
X598 2845 1 2 2678 BUF1S $T=478640 840120 1 180 $X=476160 $Y=839740
X599 2842 1 2 392 BUF1S $T=479880 739320 0 0 $X=479880 $Y=738940
X600 2866 1 2 2680 BUF1S $T=482360 840120 0 180 $X=479880 $Y=834700
X601 361 1 2 391 BUF1S $T=481120 880440 0 0 $X=481120 $Y=880060
X602 2874 1 2 2656 BUF1S $T=484220 799800 0 180 $X=481740 $Y=794380
X603 2841 1 2 2670 BUF1S $T=484220 809880 1 180 $X=481740 $Y=809500
X604 2876 1 2 2692 BUF1S $T=486080 789720 0 180 $X=483600 $Y=784300
X605 2882 1 2 394 BUF1S $T=487320 880440 0 180 $X=484840 $Y=875020
X606 2882 1 2 2717 BUF1S $T=489180 870360 1 180 $X=486700 $Y=869980
X607 2902 1 2 2842 BUF1S $T=490420 769560 1 0 $X=490420 $Y=764140
X608 2824 1 2 2923 BUF1S $T=492900 870360 0 0 $X=492900 $Y=869980
X609 403 1 2 344 BUF1S $T=494140 900600 1 0 $X=494140 $Y=895180
X610 2956 1 2 2684 BUF1S $T=502200 870360 1 180 $X=499720 $Y=869980
X611 2580 1 2 2952 BUF1S $T=500340 809880 0 0 $X=500340 $Y=809500
X612 2965 1 2 2845 BUF1S $T=502820 830040 1 180 $X=500340 $Y=829660
X613 2828 1 2 2966 BUF1S $T=500960 860280 1 0 $X=500960 $Y=854860
X614 2937 1 2 2874 BUF1S $T=503440 809880 1 0 $X=503440 $Y=804460
X615 2999 1 2 2956 BUF1S $T=507160 880440 0 180 $X=504680 $Y=875020
X616 3004 1 2 2841 BUF1S $T=509020 809880 0 180 $X=506540 $Y=804460
X617 2242 1 2 426 BUF1S $T=507160 749400 0 0 $X=507160 $Y=749020
X618 3003 1 2 404 BUF1S $T=509020 880440 0 0 $X=509020 $Y=880060
X619 2977 1 2 2876 BUF1S $T=512120 789720 0 180 $X=509640 $Y=784300
X620 2907 1 2 371 BUF1S $T=512740 890520 0 180 $X=510260 $Y=885100
X621 3010 1 2 2986 BUF1S $T=512120 759480 0 0 $X=512120 $Y=759100
X622 3035 1 2 2951 BUF1S $T=515220 769560 0 180 $X=512740 $Y=764140
X623 2907 1 2 431 BUF1S $T=513360 890520 1 0 $X=513360 $Y=885100
X624 2902 1 2 3010 BUF1S $T=513980 779640 1 0 $X=513980 $Y=774220
X625 429 1 2 3021 BUF1S $T=513980 840120 1 0 $X=513980 $Y=834700
X626 3061 1 2 2867 BUF1S $T=520180 779640 0 180 $X=517700 $Y=774220
X627 3068 1 2 2773 BUF1S $T=521420 850200 1 180 $X=518940 $Y=849820
X628 433 1 2 2993 BUF1S $T=520800 789720 1 0 $X=520800 $Y=784300
X629 2929 1 2 3054 BUF1S $T=520800 799800 0 0 $X=520800 $Y=799420
X630 3068 1 2 380 BUF1S $T=523280 880440 1 180 $X=520800 $Y=880060
X631 3093 1 2 2866 BUF1S $T=525140 830040 0 180 $X=522660 $Y=824620
X632 3094 1 2 2871 BUF1S $T=525140 840120 1 180 $X=522660 $Y=839740
X633 2895 1 2 3053 BUF1S $T=528240 840120 0 0 $X=528240 $Y=839740
X634 3010 1 2 3135 BUF1S $T=529480 779640 0 0 $X=529480 $Y=779260
X635 2947 1 2 3157 BUF1S $T=535060 819960 1 0 $X=535060 $Y=814540
X636 3092 1 2 447 BUF1S $T=537540 870360 0 180 $X=535060 $Y=864940
X637 3177 1 2 449 BUF1S $T=539400 840120 1 180 $X=536920 $Y=839740
X638 3176 1 2 3148 BUF1S $T=538780 779640 1 0 $X=538780 $Y=774220
X639 3161 1 2 3092 BUF1S $T=542500 809880 1 0 $X=542500 $Y=804460
X640 3204 1 2 3074 BUF1S $T=546220 749400 1 180 $X=543740 $Y=749020
X641 3208 1 2 452 BUF1S $T=548080 850200 1 180 $X=545600 $Y=849820
X642 3227 1 2 3141 BUF1S $T=551180 850200 1 180 $X=548700 $Y=849820
X643 3252 1 2 3109 BUF1S $T=555520 739320 0 180 $X=553040 $Y=733900
X644 3250 1 2 446 BUF1S $T=555520 890520 0 180 $X=553040 $Y=885100
X645 3256 1 2 3061 BUF1S $T=557380 779640 1 180 $X=554900 $Y=779260
X646 3196 1 2 3227 BUF1S $T=556140 830040 0 0 $X=556140 $Y=829660
X647 3199 1 2 3283 BUF1S $T=559240 799800 1 0 $X=559240 $Y=794380
X648 3271 1 2 480 BUF1S $T=559240 890520 0 0 $X=559240 $Y=890140
X649 3287 1 2 3215 BUF1S $T=562340 840120 0 180 $X=559860 $Y=834700
X650 475 1 2 454 BUF1S $T=562340 819960 1 0 $X=562340 $Y=814540
X651 3287 1 2 3271 BUF1S $T=566060 860280 1 180 $X=563580 $Y=859900
X652 3214 1 2 3270 BUF1S $T=565440 870360 1 0 $X=565440 $Y=864940
X653 488 1 2 3280 BUF1S $T=566060 819960 1 0 $X=566060 $Y=814540
X654 3190 1 2 3332 BUF1S $T=568540 799800 1 0 $X=568540 $Y=794380
X655 3297 1 2 493 BUF1S $T=568540 890520 0 0 $X=568540 $Y=890140
X656 3291 1 2 3350 BUF1S $T=572260 870360 0 0 $X=572260 $Y=869980
X657 3352 1 2 3317 BUF1S $T=573500 840120 0 0 $X=573500 $Y=839740
X658 3003 1 2 507 BUF1S $T=574120 799800 0 0 $X=574120 $Y=799420
X659 3370 1 2 3345 BUF1S $T=577220 870360 1 180 $X=574740 $Y=869980
X660 3370 1 2 511 BUF1S $T=579080 870360 0 0 $X=579080 $Y=869980
X661 3283 1 2 3419 BUF1S $T=586520 799800 0 180 $X=584040 $Y=794380
X662 3389 1 2 3452 BUF1S $T=590860 769560 0 0 $X=590860 $Y=769180
X663 494 1 2 3408 BUF1S $T=590860 819960 1 0 $X=590860 $Y=814540
X664 3385 1 2 3458 BUF1S $T=592100 819960 0 0 $X=592100 $Y=819580
X665 3225 1 2 3473 BUF1S $T=594580 809880 1 0 $X=594580 $Y=804460
X666 540 1 2 3475 BUF1S $T=595200 840120 1 0 $X=595200 $Y=834700
X667 3490 1 2 3204 BUF1S $T=598920 769560 0 180 $X=596440 $Y=764140
X668 3484 1 2 3432 BUF1S $T=598920 850200 1 180 $X=596440 $Y=849820
X669 519 1 2 520 BUF1S $T=597060 809880 1 0 $X=597060 $Y=804460
X670 3472 1 2 3461 BUF1S $T=597680 890520 0 0 $X=597680 $Y=890140
X671 3484 1 2 538 BUF1S $T=598920 870360 0 0 $X=598920 $Y=869980
X672 3250 1 2 551 BUF1S $T=600160 799800 1 0 $X=600160 $Y=794380
X673 3472 1 2 500 BUF1S $T=604500 779640 1 0 $X=604500 $Y=774220
X674 3428 1 2 3501 BUF1S $T=605120 860280 0 0 $X=605120 $Y=859900
X675 3485 1 2 3464 BUF1S $T=610700 860280 0 180 $X=608220 $Y=854860
X676 3528 1 2 3584 BUF1S $T=616900 799800 1 0 $X=616900 $Y=794380
X677 3473 1 2 3582 BUF1S $T=618760 880440 0 0 $X=618760 $Y=880060
X678 3606 1 2 3527 BUF1S $T=623100 739320 1 180 $X=620620 $Y=738940
X679 577 1 2 562 BUF1S $T=624960 900600 0 180 $X=622480 $Y=895180
X680 3463 1 2 589 BUF1S $T=624960 749400 0 0 $X=624960 $Y=749020
X681 590 1 2 3482 BUF1S $T=627440 749400 0 0 $X=627440 $Y=749020
X682 2949 1 2 3566 BUF1S $T=629920 870360 0 180 $X=627440 $Y=864940
X683 3658 1 2 3638 BUF1S $T=630540 860280 1 0 $X=630540 $Y=854860
X684 3467 1 2 607 BUF1S $T=633020 850200 1 0 $X=633020 $Y=844780
X685 603 1 2 593 BUF1S $T=635500 860280 0 180 $X=633020 $Y=854860
X686 3664 1 2 604 BUF1S $T=633020 870360 0 0 $X=633020 $Y=869980
X687 3555 1 2 3654 BUF1S $T=636120 819960 0 0 $X=636120 $Y=819580
X688 3679 1 2 3647 BUF1S $T=637360 799800 0 0 $X=637360 $Y=799420
X689 3662 1 2 3554 BUF1S $T=637980 749400 0 0 $X=637980 $Y=749020
X690 3678 1 2 3563 BUF1S $T=640460 779640 1 180 $X=637980 $Y=779260
X691 3706 1 2 3528 BUF1S $T=642940 789720 1 180 $X=640460 $Y=789340
X692 3735 1 2 3577 BUF1S $T=649140 759480 0 180 $X=646660 $Y=754060
X693 3393 1 2 3714 BUF1S $T=646660 789720 0 0 $X=646660 $Y=789340
X694 3693 1 2 3549 BUF1S $T=649760 799800 0 180 $X=647280 $Y=794380
X695 3712 1 2 3644 BUF1S $T=649140 779640 1 0 $X=649140 $Y=774220
X696 3746 1 2 569 BUF1S $T=652240 729240 1 180 $X=649760 $Y=728860
X697 639 1 2 3713 BUF1S $T=652240 729240 0 0 $X=652240 $Y=728860
X698 3773 1 2 3767 BUF1S $T=658440 840120 0 180 $X=655960 $Y=834700
X699 3729 1 2 637 BUF1S $T=658440 880440 0 180 $X=655960 $Y=875020
X700 3800 1 2 3712 BUF1S $T=663400 779640 1 180 $X=660920 $Y=779260
X701 654 1 2 3764 BUF1S $T=663400 830040 0 180 $X=660920 $Y=824620
X702 3822 1 2 3606 BUF1S $T=665260 739320 1 180 $X=662780 $Y=738940
X703 3828 1 2 3693 BUF1S $T=665260 799800 0 180 $X=662780 $Y=794380
X704 3794 1 2 651 BUF1S $T=666500 729240 0 0 $X=666500 $Y=728860
X705 3679 1 2 3832 BUF1S $T=666500 789720 0 0 $X=666500 $Y=789340
X706 3825 1 2 3808 BUF1S $T=668360 870360 1 0 $X=668360 $Y=864940
X707 666 1 2 3837 BUF1S $T=668360 890520 1 0 $X=668360 $Y=885100
X708 3842 1 2 3608 BUF1S $T=672700 769560 1 180 $X=670220 $Y=769180
X709 3867 1 2 3678 BUF1S $T=675180 769560 1 180 $X=672700 $Y=769180
X710 685 1 2 605 BUF1S $T=677660 729240 0 180 $X=675180 $Y=723820
X711 3794 1 2 3829 BUF1S $T=675180 759480 0 0 $X=675180 $Y=759100
X712 3906 1 2 3662 BUF1S $T=679520 749400 0 180 $X=677040 $Y=743980
X713 3748 1 2 3888 BUF1S $T=677660 799800 1 0 $X=677660 $Y=794380
X714 3887 1 2 3797 BUF1S $T=678280 819960 1 0 $X=678280 $Y=814540
X715 3887 1 2 3750 BUF1S $T=681380 809880 1 180 $X=678900 $Y=809500
X716 3896 1 2 3921 BUF1S $T=682620 860280 1 0 $X=682620 $Y=854860
X717 690 1 2 3896 BUF1S $T=685720 890520 1 180 $X=683240 $Y=890140
X718 3903 1 2 3935 BUF1S $T=686960 860280 1 0 $X=686960 $Y=854860
X719 3947 1 2 3706 BUF1S $T=691920 769560 1 180 $X=689440 $Y=769180
X720 3955 1 2 3951 BUF1S $T=690060 850200 1 0 $X=690060 $Y=844780
X721 3896 1 2 3898 BUF1S $T=691300 819960 1 0 $X=691300 $Y=814540
X722 3797 1 2 3955 BUF1S $T=695020 819960 1 0 $X=695020 $Y=814540
X723 426 1 2 3910 BUF1S $T=695640 759480 0 0 $X=695640 $Y=759100
X724 3955 1 2 4007 BUF1S $T=697500 809880 0 0 $X=697500 $Y=809500
X725 4027 1 2 3739 BUF1S $T=702460 749400 1 180 $X=699980 $Y=749020
X726 4034 1 2 3894 BUF1S $T=702460 759480 0 180 $X=699980 $Y=754060
X727 4039 1 2 3735 BUF1S $T=704940 749400 1 180 $X=702460 $Y=749020
X728 4050 1 2 722 BUF1S $T=708660 880440 1 0 $X=708660 $Y=875020
X729 4088 1 2 3173 BUF1S $T=712380 870360 1 180 $X=709900 $Y=869980
X730 4050 1 2 4009 BUF1S $T=712380 860280 1 0 $X=712380 $Y=854860
X731 748 1 2 671 BUF1S $T=716100 870360 0 180 $X=713620 $Y=864940
X732 749 1 2 655 BUF1S $T=716720 870360 1 180 $X=714240 $Y=869980
X733 4118 1 2 4027 BUF1S $T=716100 789720 1 0 $X=716100 $Y=784300
X734 4007 1 2 4129 BUF1S $T=717960 789720 0 0 $X=717960 $Y=789340
X735 4007 1 2 4139 BUF1S $T=721060 809880 0 0 $X=721060 $Y=809500
X736 3609 1 2 4144 BUF1S $T=722300 830040 0 0 $X=722300 $Y=829660
X737 762 1 2 768 BUF1S $T=723540 729240 1 0 $X=723540 $Y=723820
X738 4162 1 2 3234 BUF1S $T=727260 749400 1 180 $X=724780 $Y=749020
X739 4159 1 2 754 BUF1S $T=727260 880440 0 180 $X=724780 $Y=875020
X740 765 1 2 3414 BUF1S $T=725400 789720 1 0 $X=725400 $Y=784300
X741 772 1 2 3333 BUF1S $T=729120 860280 1 180 $X=726640 $Y=859900
X742 4127 1 2 4159 BUF1S $T=730980 840120 1 180 $X=728500 $Y=839740
X743 4179 1 2 3941 BUF1S $T=732220 799800 0 180 $X=729740 $Y=794380
X744 4176 1 2 4180 BUF1S $T=729740 840120 1 0 $X=729740 $Y=834700
X745 4139 1 2 4193 BUF1S $T=730360 799800 0 0 $X=730360 $Y=799420
X746 4184 1 2 4197 BUF1S $T=731600 860280 1 0 $X=731600 $Y=854860
X747 4199 1 2 4012 BUF1S $T=734700 799800 0 180 $X=732220 $Y=794380
X748 4139 1 2 4192 BUF1S $T=732220 819960 0 0 $X=732220 $Y=819580
X749 795 1 2 4201 BUF1S $T=739660 739320 0 180 $X=737180 $Y=733900
X750 4264 1 2 778 BUF1S $T=747100 880440 0 180 $X=744620 $Y=875020
X751 2949 1 2 4198 BUF1S $T=745860 870360 1 0 $X=745860 $Y=864940
X752 4234 1 2 4264 BUF1S $T=748340 830040 0 0 $X=748340 $Y=829660
X753 827 1 2 4088 BUF1S $T=752680 860280 0 180 $X=750200 $Y=854860
X754 4312 1 2 3177 BUF1S $T=755160 799800 1 180 $X=752680 $Y=799420
X755 4174 1 2 828 BUF1S $T=753920 840120 1 0 $X=753920 $Y=834700
X756 4307 1 2 832 BUF1S $T=754540 729240 0 0 $X=754540 $Y=728860
X757 4317 1 2 4123 BUF1S $T=761980 880440 0 180 $X=759500 $Y=875020
X758 822 1 2 4317 BUF1S $T=764460 890520 0 180 $X=761980 $Y=885100
X759 4334 1 2 4326 BUF1S $T=764460 749400 0 0 $X=764460 $Y=749020
X760 4317 1 2 4330 BUF1S $T=764460 870360 0 0 $X=764460 $Y=869980
X761 4359 1 2 838 BUF1S $T=764460 890520 0 0 $X=764460 $Y=890140
X762 4330 1 2 4304 BUF1S $T=767560 850200 0 180 $X=765080 $Y=844780
X763 4304 1 2 4382 BUF1S $T=766320 830040 0 0 $X=766320 $Y=829660
X764 4391 1 2 4407 BUF1S $T=771280 809880 1 0 $X=771280 $Y=804460
X765 4343 1 2 4337 BUF1S $T=773140 890520 1 0 $X=773140 $Y=885100
X766 3208 1 2 868 BUF1S $T=777480 850200 1 180 $X=775000 $Y=849820
X767 857 1 2 4412 BUF1S $T=775620 789720 0 0 $X=775620 $Y=789340
X768 4224 1 2 4467 BUF1S $T=783680 779640 0 0 $X=783680 $Y=779260
X769 4467 1 2 4433 BUF1S $T=786780 769560 1 0 $X=786780 $Y=764140
X770 4243 1 2 878 BUF1S $T=788020 890520 0 0 $X=788020 $Y=890140
X771 4448 1 2 4539 BUF1S $T=792360 789720 1 0 $X=792360 $Y=784300
X772 4482 1 2 4425 BUF1S $T=792360 870360 0 0 $X=792360 $Y=869980
X773 4512 1 2 903 BUF1S $T=792360 890520 1 0 $X=792360 $Y=885100
X774 4474 1 2 4540 BUF1S $T=794840 860280 0 0 $X=794840 $Y=859900
X775 4491 1 2 904 BUF1S $T=794840 900600 1 0 $X=794840 $Y=895180
X776 4487 1 2 4498 BUF1S $T=798560 789720 1 180 $X=796080 $Y=789340
X777 4467 1 2 4576 BUF1S $T=797940 779640 1 0 $X=797940 $Y=774220
X778 4585 1 2 4455 BUF1S $T=801040 749400 1 180 $X=798560 $Y=749020
X779 4583 1 2 4462 BUF1S $T=801660 830040 1 180 $X=799180 $Y=829660
X780 4422 1 2 4575 BUF1S $T=799800 759480 0 0 $X=799800 $Y=759100
X781 4608 1 2 4560 BUF1S $T=805380 789720 1 180 $X=802900 $Y=789340
X782 4480 1 2 4646 BUF1S $T=807860 860280 0 0 $X=807860 $Y=859900
X783 4576 1 2 4639 BUF1S $T=810340 779640 1 0 $X=810340 $Y=774220
X784 4556 1 2 4461 BUF1S $T=810960 880440 0 0 $X=810960 $Y=880060
X785 776 1 2 4655 BUF1S $T=812200 779640 0 0 $X=812200 $Y=779260
X786 4510 1 2 4636 BUF1S $T=812200 799800 1 0 $X=812200 $Y=794380
X787 4574 1 2 4668 BUF1S $T=814060 739320 1 0 $X=814060 $Y=733900
X788 458 1 2 4681 BUF1S $T=814060 850200 0 0 $X=814060 $Y=849820
X789 4381 1 2 4687 BUF1S $T=815920 799800 1 0 $X=815920 $Y=794380
X790 4688 1 2 4583 BUF1S $T=818400 819960 1 180 $X=815920 $Y=819580
X791 4688 1 2 4582 BUF1S $T=818400 830040 0 180 $X=815920 $Y=824620
X792 887 1 2 938 BUF1S $T=816540 900600 1 0 $X=816540 $Y=895180
X793 935 1 2 939 BUF1S $T=817160 729240 0 0 $X=817160 $Y=728860
X794 4699 1 2 4566 BUF1S $T=820260 749400 0 180 $X=817780 $Y=743980
X795 940 1 2 4708 BUF1S $T=819020 900600 1 0 $X=819020 $Y=895180
X796 4705 1 2 4649 BUF1S $T=821500 860280 1 0 $X=821500 $Y=854860
X797 4716 1 2 4702 BUF1S $T=824600 870360 1 0 $X=824600 $Y=864940
X798 4730 1 2 4692 BUF1S $T=825840 850200 0 0 $X=825840 $Y=849820
X799 4712 1 2 4688 BUF1S $T=837000 850200 1 180 $X=834520 $Y=849820
X800 4608 1 2 4801 BUF1S $T=835140 789720 1 0 $X=835140 $Y=784300
X801 4740 1 2 4717 BUF1S $T=835140 799800 0 0 $X=835140 $Y=799420
X802 4645 1 2 960 BUF1S $T=837000 729240 0 0 $X=837000 $Y=728860
X803 765 1 2 957 BUF1S $T=837000 779640 1 0 $X=837000 $Y=774220
X804 4763 1 2 961 BUF1S $T=837620 880440 1 0 $X=837620 $Y=875020
X805 4699 1 2 964 BUF1S $T=838860 739320 1 0 $X=838860 $Y=733900
X806 4539 1 2 4820 BUF1S $T=838860 789720 1 0 $X=838860 $Y=784300
X807 4662 1 2 965 BUF1S $T=838860 799800 0 0 $X=838860 $Y=799420
X808 4821 1 2 4450 BUF1S $T=841340 819960 0 180 $X=838860 $Y=814540
X809 4407 1 2 4837 BUF1S $T=838860 819960 0 0 $X=838860 $Y=819580
X810 4731 1 2 4788 BUF1S $T=843200 860280 1 180 $X=840720 $Y=859900
X811 4716 1 2 4830 BUF1S $T=840720 870360 0 0 $X=840720 $Y=869980
X812 4825 1 2 4857 BUF1S $T=845680 870360 1 0 $X=845680 $Y=864940
X813 4721 1 2 4893 BUF1S $T=849400 759480 0 0 $X=849400 $Y=759100
X814 4585 1 2 4887 BUF1S $T=851260 749400 0 0 $X=851260 $Y=749020
X815 4725 1 2 4847 BUF1S $T=851260 769560 1 0 $X=851260 $Y=764140
X816 4814 1 2 4897 BUF1S $T=852500 850200 1 0 $X=852500 $Y=844780
X817 4700 1 2 4890 BUF1S $T=853120 739320 1 0 $X=853120 $Y=733900
X818 4575 1 2 4903 BUF1S $T=853120 759480 0 0 $X=853120 $Y=759100
X819 4899 1 2 4888 BUF1S $T=854980 749400 0 0 $X=854980 $Y=749020
X820 4720 1 2 4908 BUF1S $T=854980 769560 1 0 $X=854980 $Y=764140
X821 4822 1 2 4910 BUF1S $T=854980 870360 0 0 $X=854980 $Y=869980
X822 4822 1 2 4882 BUF1S $T=854980 880440 1 0 $X=854980 $Y=875020
X823 4835 1 2 4870 BUF1S $T=855600 900600 1 0 $X=855600 $Y=895180
X824 4720 1 2 4915 BUF1S $T=856220 840120 1 0 $X=856220 $Y=834700
X825 4731 1 2 4916 BUF1S $T=856220 860280 0 0 $X=856220 $Y=859900
X826 4918 1 2 4849 BUF1S $T=859320 739320 0 180 $X=856840 $Y=733900
X827 4919 1 2 4741 BUF1S $T=859320 819960 0 180 $X=856840 $Y=814540
X828 4839 1 2 4919 BUF1S $T=856840 840120 0 0 $X=856840 $Y=839740
X829 4831 1 2 4945 BUF1S $T=863040 880440 1 0 $X=863040 $Y=875020
X830 4919 1 2 4900 BUF1S $T=863660 819960 1 0 $X=863660 $Y=814540
X831 4933 1 2 4960 BUF1S $T=864900 799800 0 0 $X=864900 $Y=799420
X832 4847 1 2 4948 BUF1S $T=865520 769560 1 0 $X=865520 $Y=764140
X833 980 1 2 4911 BUF1S $T=866760 890520 1 0 $X=866760 $Y=885100
X834 4824 1 2 4982 BUF1S $T=867380 870360 1 0 $X=867380 $Y=864940
X835 4972 1 2 4983 BUF1S $T=869240 749400 1 0 $X=869240 $Y=743980
X836 980 1 2 990 BUF1S $T=869240 890520 1 0 $X=869240 $Y=885100
X837 4800 1 2 4981 BUF1S $T=872340 850200 1 0 $X=872340 $Y=844780
X838 980 1 2 972 BUF1S $T=877300 890520 0 0 $X=877300 $Y=890140
X839 4900 1 2 5020 BUF1S $T=877920 809880 1 0 $X=877920 $Y=804460
X840 4911 1 2 4927 BUF1S $T=881020 880440 0 180 $X=878540 $Y=875020
X841 4927 1 2 5021 BUF1S $T=880400 850200 0 0 $X=880400 $Y=849820
X842 5121 1 2 5061 BUF1S $T=895280 830040 1 0 $X=895280 $Y=824620
X843 4911 1 2 5101 BUF1S $T=895280 880440 1 0 $X=895280 $Y=875020
X844 5021 1 2 5117 BUF1S $T=897760 830040 1 0 $X=897760 $Y=824620
X845 5144 1 2 5150 BUF1S $T=899000 830040 0 0 $X=899000 $Y=829660
X846 5147 1 2 5169 BUF1S $T=902100 870360 1 0 $X=902100 $Y=864940
X847 1018 1 2 5008 BUF1S $T=905820 789720 0 180 $X=903340 $Y=784300
X848 5185 1 2 5016 BUF1S $T=907060 840120 0 180 $X=904580 $Y=834700
X849 5183 1 2 5095 BUF1S $T=908300 860280 0 180 $X=905820 $Y=854860
X850 5042 1 2 5034 BUF1S $T=908920 769560 0 180 $X=906440 $Y=764140
X851 4953 1 2 5195 BUF1S $T=906440 789720 1 0 $X=906440 $Y=784300
X852 5181 1 2 5042 BUF1S $T=911400 789720 0 180 $X=908920 $Y=784300
X853 5185 1 2 991 BUF1S $T=911400 840120 0 0 $X=911400 $Y=839740
X854 5162 1 2 1042 BUF1S $T=913880 830040 1 0 $X=913880 $Y=824620
X855 5117 1 2 5226 BUF1S $T=915120 830040 0 0 $X=915120 $Y=829660
X856 5225 1 2 1036 BUF1S $T=916980 739320 1 0 $X=916980 $Y=733900
X857 5253 1 2 5225 BUF1S $T=923180 779640 0 180 $X=920700 $Y=774220
X858 5227 1 2 5194 BUF1S $T=920700 860280 1 0 $X=920700 $Y=854860
X859 5101 1 2 5227 BUF1S $T=923180 860280 1 180 $X=920700 $Y=859900
X860 5241 1 2 5274 BUF1S $T=927520 759480 1 0 $X=927520 $Y=754060
X861 5225 1 2 5294 BUF1S $T=928760 749400 0 0 $X=928760 $Y=749020
X862 5269 1 2 5304 BUF1S $T=929380 870360 1 0 $X=929380 $Y=864940
X863 1053 1 2 5261 BUF1S $T=933720 900600 0 180 $X=931240 $Y=895180
X864 5179 1 2 1054 BUF1S $T=933100 739320 0 0 $X=933100 $Y=738940
X865 5233 1 2 5330 BUF1S $T=933100 779640 0 0 $X=933100 $Y=779260
X866 5269 1 2 5323 BUF1S $T=933720 860280 1 0 $X=933720 $Y=854860
X867 5242 1 2 5337 BUF1S $T=934340 830040 1 0 $X=934340 $Y=824620
X868 5233 1 2 1055 BUF1S $T=934960 729240 1 0 $X=934960 $Y=723820
X869 5212 1 2 5338 BUF1S $T=934960 759480 1 0 $X=934960 $Y=754060
X870 5266 1 2 1057 BUF1S $T=934960 890520 0 0 $X=934960 $Y=890140
X871 5212 1 2 5345 BUF1S $T=936200 769560 1 0 $X=936200 $Y=764140
X872 5266 1 2 5291 BUF1S $T=936200 860280 1 0 $X=936200 $Y=854860
X873 5350 1 2 5367 BUF1S $T=938680 870360 1 0 $X=938680 $Y=864940
X874 5360 1 2 5381 BUF1S $T=939920 850200 1 0 $X=939920 $Y=844780
X875 5309 1 2 5355 BUF1S $T=945500 759480 1 0 $X=945500 $Y=754060
X876 5337 1 2 5361 BUF1S $T=945500 799800 0 0 $X=945500 $Y=799420
X877 5267 1 2 5427 BUF1S $T=947360 779640 1 0 $X=947360 $Y=774220
X878 4976 1 2 1074 BUF1S $T=948600 809880 1 0 $X=948600 $Y=804460
X879 5434 1 2 1075 BUF1S $T=951080 890520 1 0 $X=951080 $Y=885100
X880 5295 1 2 5461 BUF1S $T=954180 739320 0 0 $X=954180 $Y=738940
X881 5453 1 2 5462 BUF1S $T=954180 779640 1 0 $X=954180 $Y=774220
X882 1078 1 2 5332 BUF1S $T=954180 880440 1 0 $X=954180 $Y=875020
X883 1082 1 2 5468 BUF1S $T=959140 870360 0 180 $X=956660 $Y=864940
X884 5326 1 2 5475 BUF1S $T=957900 759480 1 0 $X=957900 $Y=754060
X885 5468 1 2 5324 BUF1S $T=961620 870360 1 180 $X=959140 $Y=869980
X886 1067 1 2 5437 BUF1S $T=963480 850200 0 180 $X=961000 $Y=844780
X887 5501 1 2 5496 BUF1S $T=961620 860280 0 0 $X=961620 $Y=859900
X888 5329 1 2 5459 BUF1S $T=962240 809880 0 0 $X=962240 $Y=809500
X889 5337 1 2 5454 BUF1S $T=963480 819960 1 0 $X=963480 $Y=814540
X890 1085 1 2 5501 BUF1S $T=964100 880440 1 0 $X=964100 $Y=875020
X891 5319 1 2 5445 BUF1S $T=964720 830040 0 0 $X=964720 $Y=829660
X892 1067 1 2 1051 BUF1S $T=964720 860280 1 0 $X=964720 $Y=854860
X893 5503 1 2 5398 BUF1S $T=967820 850200 0 0 $X=967820 $Y=849820
X894 5294 1 2 5568 BUF1S $T=972160 739320 0 0 $X=972160 $Y=738940
X895 1097 1 2 5557 BUF1S $T=974640 779640 1 180 $X=972160 $Y=779260
X896 1070 1 2 5536 BUF1S $T=974020 900600 1 0 $X=974020 $Y=895180
X897 5580 1 2 5587 BUF1S $T=974640 769560 1 0 $X=974640 $Y=764140
X898 1080 1 2 5600 BUF1S $T=975880 749400 1 0 $X=975880 $Y=743980
X899 5582 1 2 5602 BUF1S $T=976500 890520 1 0 $X=976500 $Y=885100
X900 5454 1 2 5608 BUF1S $T=977740 799800 0 0 $X=977740 $Y=799420
X901 1098 1 2 5497 BUF1S $T=985180 769560 1 180 $X=982700 $Y=769180
X902 5639 1 2 5460 BUF1S $T=987040 840120 0 180 $X=984560 $Y=834700
X903 5647 1 2 5648 BUF1S $T=988900 809880 0 0 $X=988900 $Y=809500
X904 5652 1 2 5661 BUF1S $T=991380 789720 0 0 $X=991380 $Y=789340
X905 4312 1 2 1113 BUF1S $T=997580 819960 1 180 $X=995100 $Y=819580
X906 5651 1 2 5639 BUF1S $T=997580 840120 0 180 $X=995100 $Y=834700
X907 892 1 2 1117 BUF1S $T=996960 830040 1 0 $X=996960 $Y=824620
X908 5701 1 2 5653 BUF1S $T=1000680 809880 0 0 $X=1000680 $Y=809500
X909 5677 1 2 5736 BUF1S $T=1001920 739320 1 0 $X=1001920 $Y=733900
X910 5719 1 2 5734 BUF1S $T=1002540 870360 1 0 $X=1002540 $Y=864940
X911 5650 1 2 5750 BUF1S $T=1004400 759480 0 0 $X=1004400 $Y=759100
X912 5755 1 2 5745 BUF1S $T=1006880 809880 0 0 $X=1006880 $Y=809500
X913 1108 1 2 5774 BUF1S $T=1007500 890520 0 0 $X=1007500 $Y=890140
X914 5757 1 2 1141 BUF1S $T=1010600 870360 0 0 $X=1010600 $Y=869980
X915 5786 1 2 5763 BUF1S $T=1011840 860280 0 0 $X=1011840 $Y=859900
X916 5700 1 2 5796 BUF1S $T=1013080 759480 1 0 $X=1013080 $Y=754060
X917 5657 1 2 5766 BUF1S $T=1015560 840120 0 180 $X=1013080 $Y=834700
X918 5693 1 2 5754 BUF1S $T=1013700 789720 0 0 $X=1013700 $Y=789340
X919 1145 1 2 1143 BUF1S $T=1016180 900600 0 180 $X=1013700 $Y=895180
X920 5736 1 2 5803 BUF1S $T=1014940 739320 0 0 $X=1014940 $Y=738940
X921 5666 1 2 5775 BUF1S $T=1014940 880440 0 0 $X=1014940 $Y=880060
X922 5741 1 2 5798 BUF1S $T=1016180 830040 0 0 $X=1016180 $Y=829660
X923 5789 1 2 5820 BUF1S $T=1018040 739320 1 0 $X=1018040 $Y=733900
X924 5817 1 2 5760 BUF1S $T=1019280 809880 0 0 $X=1019280 $Y=809500
X925 5756 1 2 5694 BUF1S $T=1021760 840120 1 0 $X=1021760 $Y=834700
X926 5844 1 2 5836 BUF1S $T=1023620 819960 1 0 $X=1023620 $Y=814540
X927 885 1 2 1159 BUF1S $T=1023620 830040 1 0 $X=1023620 $Y=824620
X928 5720 1 2 5863 BUF1S $T=1025480 759480 1 0 $X=1025480 $Y=754060
X929 5501 1 2 1149 BUF1S $T=1025480 900600 1 0 $X=1025480 $Y=895180
X930 5796 1 2 5878 BUF1S $T=1027960 759480 1 0 $X=1027960 $Y=754060
X931 5872 1 2 5835 BUF1S $T=1027960 830040 1 0 $X=1027960 $Y=824620
X932 5733 1 2 5888 BUF1S $T=1029200 789720 1 0 $X=1029200 $Y=784300
X933 1104 1 2 1169 BUF1S $T=1030440 830040 1 0 $X=1030440 $Y=824620
X934 5879 1 2 5680 BUF1S $T=1030440 850200 0 0 $X=1030440 $Y=849820
X935 5848 1 2 5865 BUF1S $T=1031060 789720 0 0 $X=1031060 $Y=789340
X936 5701 1 2 5900 BUF1S $T=1031060 809880 1 0 $X=1031060 $Y=804460
X937 5902 1 2 5926 BUF1S $T=1032920 850200 0 0 $X=1032920 $Y=849820
X938 5914 1 2 5930 BUF1S $T=1034160 890520 0 0 $X=1034160 $Y=890140
X939 5923 1 2 1166 BUF1S $T=1040360 860280 0 180 $X=1037880 $Y=854860
X940 5926 1 2 1177 BUF1S $T=1037880 880440 1 0 $X=1037880 $Y=875020
X941 1180 1 2 5853 BUF1S $T=1042220 729240 0 180 $X=1039740 $Y=723820
X942 5943 1 2 5949 BUF1S $T=1039740 799800 1 0 $X=1039740 $Y=794380
X943 5884 1 2 5963 BUF1S $T=1040360 860280 1 0 $X=1040360 $Y=854860
X944 5949 1 2 5819 BUF1S $T=1044080 779640 0 180 $X=1041600 $Y=774220
X945 1178 1 2 5877 BUF1S $T=1042220 729240 1 0 $X=1042220 $Y=723820
X946 5925 1 2 5928 BUF1S $T=1044080 850200 0 0 $X=1044080 $Y=849820
X947 5501 1 2 5935 BUF1S $T=1045940 830040 1 0 $X=1045940 $Y=824620
X948 5981 1 2 5965 BUF1S $T=1045940 870360 0 0 $X=1045940 $Y=869980
X949 5956 1 2 1185 BUF1S $T=1046560 850200 0 0 $X=1046560 $Y=849820
X950 5911 1 2 5968 BUF1S $T=1047800 739320 0 0 $X=1047800 $Y=738940
X951 5962 1 2 5940 BUF1S $T=1048420 830040 1 0 $X=1048420 $Y=824620
X952 6003 1 2 5943 BUF1S $T=1050900 819960 0 0 $X=1050900 $Y=819580
X953 5797 1 2 6020 BUF1S $T=1052140 830040 1 0 $X=1052140 $Y=824620
X954 5802 1 2 6026 BUF1S $T=1052140 830040 0 0 $X=1052140 $Y=829660
X955 5926 1 2 6024 BUF1S $T=1052760 860280 1 0 $X=1052760 $Y=854860
X956 5949 1 2 5974 BUF1S $T=1055860 759480 1 180 $X=1053380 $Y=759100
X957 1148 1 2 5864 BUF1S $T=1056480 779640 1 180 $X=1054000 $Y=779260
X958 5967 1 2 5889 BUF1S $T=1054620 830040 1 0 $X=1054620 $Y=824620
X959 5666 1 2 6036 BUF1S $T=1055240 880440 0 0 $X=1055240 $Y=880060
X960 5794 1 2 6041 BUF1S $T=1055860 880440 1 0 $X=1055860 $Y=875020
X961 5923 1 2 6048 BUF1S $T=1057100 850200 0 0 $X=1057100 $Y=849820
X962 1162 1 2 1194 BUF1S $T=1060820 729240 1 0 $X=1060820 $Y=723820
X963 5900 1 2 6082 BUF1S $T=1063920 809880 1 0 $X=1063920 $Y=804460
X964 1148 1 2 1198 BUF1S $T=1064540 900600 1 0 $X=1064540 $Y=895180
X965 6069 1 2 6050 BUF1S $T=1065780 769560 0 0 $X=1065780 $Y=769180
X966 5863 1 2 6091 BUF1S $T=1066400 759480 1 0 $X=1066400 $Y=754060
X967 5955 1 2 6104 BUF1S $T=1067640 809880 0 0 $X=1067640 $Y=809500
X968 6033 1 2 6088 BUF1S $T=1068880 789720 0 0 $X=1068880 $Y=789340
X969 6107 1 2 6102 BUF1S $T=1073840 850200 0 0 $X=1073840 $Y=849820
X970 6090 1 2 6139 BUF1S $T=1075700 739320 1 0 $X=1075700 $Y=733900
X971 6088 1 2 6146 BUF1S $T=1086240 769560 0 180 $X=1083760 $Y=764140
X972 6123 1 2 6140 BUF1S $T=1085620 799800 0 0 $X=1085620 $Y=799420
X973 6127 1 2 6188 BUF1S $T=1085620 830040 1 0 $X=1085620 $Y=824620
X974 6206 1 2 6128 BUF1S $T=1091820 840120 1 180 $X=1089340 $Y=839740
X975 1220 1 2 6107 BUF1S $T=1092440 789720 0 0 $X=1092440 $Y=789340
X976 6088 1 2 6224 BUF1S $T=1094300 769560 1 0 $X=1094300 $Y=764140
X977 6188 1 2 6210 BUF1S $T=1099880 819960 1 0 $X=1099880 $Y=814540
X978 6223 1 2 6280 BUF1S $T=1101740 890520 1 0 $X=1101740 $Y=885100
X979 6269 1 2 6298 BUF1S $T=1104220 819960 1 0 $X=1104220 $Y=814540
X980 1241 1 2 6206 BUF1S $T=1107940 890520 1 180 $X=1105460 $Y=890140
X981 6328 1 2 6352 BUF1S $T=1114140 860280 1 0 $X=1114140 $Y=854860
X982 1247 1 2 6362 BUF1S $T=1114140 880440 1 0 $X=1114140 $Y=875020
X983 6140 1 2 6369 BUF1S $T=1116000 779640 1 0 $X=1116000 $Y=774220
X984 6362 1 2 6251 BUF1S $T=1129020 850200 0 180 $X=1126540 $Y=844780
X985 6367 1 2 6371 BUF1S $T=1126540 890520 1 0 $X=1126540 $Y=885100
X986 1331 1 2 1328 DELB $T=223200 729240 0 0 $X=223200 $Y=728860
X987 1343 1 2 1363 DELB $T=225060 739320 1 0 $X=225060 $Y=733900
X988 1375 1 2 21 DELB $T=230020 729240 0 0 $X=230020 $Y=728860
X989 1444 1 2 1441 DELB $T=240560 749400 1 0 $X=240560 $Y=743980
X990 1465 1 2 1471 DELB $T=245520 739320 1 0 $X=245520 $Y=733900
X991 1895 1 2 1919 DELB $T=321160 809880 1 0 $X=321160 $Y=804460
X992 1930 1 2 1944 DELB $T=327980 739320 0 0 $X=327980 $Y=738940
X993 1978 1 2 1961 DELB $T=344100 799800 0 0 $X=344100 $Y=799420
X994 2099 1 2 2115 DELB $T=360840 819960 0 0 $X=360840 $Y=819580
X995 2251 1 2 2275 DELB $T=375100 870360 1 0 $X=375100 $Y=864940
X996 2355 1 2 2384 DELB $T=389980 850200 1 0 $X=389980 $Y=844780
X997 264 1 2 272 DELB $T=389980 900600 1 0 $X=389980 $Y=895180
X998 2484 1 2 2519 DELB $T=411060 789720 0 0 $X=411060 $Y=789340
X999 2493 1 2 2520 DELB $T=411060 840120 1 0 $X=411060 $Y=834700
X1000 2533 1 2 2551 DELB $T=417880 870360 0 0 $X=417880 $Y=869980
X1001 2543 1 2 2558 DELB $T=419740 769560 0 0 $X=419740 $Y=769180
X1002 2549 1 2 2570 DELB $T=421600 789720 0 0 $X=421600 $Y=789340
X1003 2552 1 2 2574 DELB $T=422220 880440 0 0 $X=422220 $Y=880060
X1004 2610 1 2 2636 DELB $T=434620 860280 0 0 $X=434620 $Y=859900
X1005 2619 1 2 2644 DELB $T=437100 789720 1 0 $X=437100 $Y=784300
X1006 2642 1 2 2666 DELB $T=441440 769560 1 0 $X=441440 $Y=764140
X1007 2704 1 2 2687 DELB $T=450120 759480 0 0 $X=450120 $Y=759100
X1008 2643 1 2 2671 DELB $T=450120 789720 0 0 $X=450120 $Y=789340
X1009 2645 1 2 2672 DELB $T=450120 830040 1 0 $X=450120 $Y=824620
X1010 2721 1 2 2745 DELB $T=455080 860280 1 0 $X=455080 $Y=854860
X1011 2729 1 2 2731 DELB $T=456320 789720 0 0 $X=456320 $Y=789340
X1012 2792 1 2 2817 DELB $T=468100 729240 1 0 $X=468100 $Y=723820
X1013 2822 1 2 2846 DELB $T=473680 769560 1 0 $X=473680 $Y=764140
X1014 2827 1 2 2800 DELB $T=474920 860280 0 0 $X=474920 $Y=859900
X1015 2757 1 2 2848 DELB $T=478640 890520 1 0 $X=478640 $Y=885100
X1016 2818 1 2 2875 DELB $T=480500 769560 1 0 $X=480500 $Y=764140
X1017 2840 1 2 2863 DELB $T=482360 830040 1 0 $X=482360 $Y=824620
X1018 2850 1 2 2832 DELB $T=482360 840120 1 0 $X=482360 $Y=834700
X1019 2861 1 2 2883 DELB $T=486080 739320 0 0 $X=486080 $Y=738940
X1020 2892 1 2 2890 DELB $T=487940 819960 1 0 $X=487940 $Y=814540
X1021 2920 1 2 2921 DELB $T=494760 819960 1 0 $X=494760 $Y=814540
X1022 2928 1 2 2904 DELB $T=496620 789720 1 0 $X=496620 $Y=784300
X1023 2934 1 2 2939 DELB $T=497860 759480 0 0 $X=497860 $Y=759100
X1024 2944 1 2 2973 DELB $T=499100 860280 0 0 $X=499100 $Y=859900
X1025 406 1 2 2953 DELB $T=499720 739320 1 0 $X=499720 $Y=733900
X1026 2954 1 2 2972 DELB $T=503440 789720 1 0 $X=503440 $Y=784300
X1027 2981 1 2 2982 DELB $T=504680 759480 0 0 $X=504680 $Y=759100
X1028 417 1 2 425 DELB $T=505300 890520 1 0 $X=505300 $Y=885100
X1029 2988 1 2 3000 DELB $T=507160 819960 0 0 $X=507160 $Y=819580
X1030 3001 1 2 2950 DELB $T=507780 850200 1 0 $X=507780 $Y=844780
X1031 3037 1 2 3038 DELB $T=514600 819960 1 0 $X=514600 $Y=814540
X1032 3031 1 2 3011 DELB $T=515220 880440 1 0 $X=515220 $Y=875020
X1033 3013 1 2 3030 DELB $T=515840 900600 1 0 $X=515840 $Y=895180
X1034 2992 1 2 3090 DELB $T=516460 840120 1 0 $X=516460 $Y=834700
X1035 3059 1 2 3085 DELB $T=519560 759480 1 0 $X=519560 $Y=754060
X1036 3078 1 2 3130 DELB $T=522660 880440 1 0 $X=522660 $Y=875020
X1037 3088 1 2 3117 DELB $T=523900 809880 1 0 $X=523900 $Y=804460
X1038 3105 1 2 3104 DELB $T=526380 830040 1 0 $X=526380 $Y=824620
X1039 3126 1 2 3125 DELB $T=529480 860280 0 0 $X=529480 $Y=859900
X1040 3129 1 2 3162 DELB $T=531960 840120 0 0 $X=531960 $Y=839740
X1041 3121 1 2 3142 DELB $T=535680 890520 0 0 $X=535680 $Y=890140
X1042 3170 1 2 3183 DELB $T=540640 729240 0 0 $X=540640 $Y=728860
X1043 3182 1 2 3205 DELB $T=541260 799800 0 0 $X=541260 $Y=799420
X1044 3206 1 2 3224 DELB $T=546220 799800 1 0 $X=546220 $Y=794380
X1045 463 1 2 467 DELB $T=548080 890520 1 0 $X=548080 $Y=885100
X1046 445 1 2 3134 DELB $T=548700 729240 0 0 $X=548700 $Y=728860
X1047 3276 1 2 3258 DELB $T=559860 759480 0 0 $X=559860 $Y=759100
X1048 478 1 2 485 DELB $T=560480 729240 1 0 $X=560480 $Y=723820
X1049 3242 1 2 3282 DELB $T=565440 880440 0 0 $X=565440 $Y=880060
X1050 3313 1 2 3337 DELB $T=566680 729240 0 0 $X=566680 $Y=728860
X1051 3289 1 2 3294 DELB $T=567920 860280 0 0 $X=567920 $Y=859900
X1052 3279 1 2 3307 DELB $T=571020 759480 1 0 $X=571020 $Y=754060
X1053 3355 1 2 3325 DELB $T=575980 759480 0 0 $X=575980 $Y=759100
X1054 505 1 2 516 DELB $T=576600 729240 1 0 $X=576600 $Y=723820
X1055 3398 1 2 3400 DELB $T=579700 809880 1 0 $X=579700 $Y=804460
X1056 3381 1 2 3391 DELB $T=582180 759480 1 0 $X=582180 $Y=754060
X1057 3402 1 2 3427 DELB $T=582180 830040 0 0 $X=582180 $Y=829660
X1058 3392 1 2 3446 DELB $T=587140 729240 0 0 $X=587140 $Y=728860
X1059 3336 1 2 3293 DELB $T=587140 870360 1 0 $X=587140 $Y=864940
X1060 531 1 2 3447 DELB $T=587760 789720 0 0 $X=587760 $Y=789340
X1061 3364 1 2 3383 DELB $T=592100 789720 1 0 $X=592100 $Y=784300
X1062 3433 1 2 3477 DELB $T=592720 870360 1 0 $X=592720 $Y=864940
X1063 3456 1 2 3481 DELB $T=593340 880440 0 0 $X=593340 $Y=880060
X1064 3500 1 2 3529 DELB $T=600780 799800 0 0 $X=600780 $Y=799420
X1065 3513 1 2 3523 DELB $T=602640 739320 0 0 $X=602640 $Y=738940
X1066 3492 1 2 3509 DELB $T=602640 789720 1 0 $X=602640 $Y=784300
X1067 3559 1 2 3580 DELB $T=613180 789720 1 0 $X=613180 $Y=784300
X1068 3560 1 2 3581 DELB $T=613180 840120 0 0 $X=613180 $Y=839740
X1069 3568 1 2 3567 DELB $T=615040 749400 0 0 $X=615040 $Y=749020
X1070 3564 1 2 3551 DELB $T=618760 759480 0 0 $X=618760 $Y=759100
X1071 3517 1 2 3595 DELB $T=620000 890520 0 0 $X=620000 $Y=890140
X1072 3689 1 2 3688 DELB $T=637360 890520 0 0 $X=637360 $Y=890140
X1073 3624 1 2 3650 DELB $T=638600 819960 0 0 $X=638600 $Y=819580
X1074 3726 1 2 3745 DELB $T=646660 890520 1 0 $X=646660 $Y=885100
X1075 3727 1 2 3732 DELB $T=647280 759480 0 0 $X=647280 $Y=759100
X1076 641 1 2 649 DELB $T=652860 900600 1 0 $X=652860 $Y=895180
X1077 3723 1 2 3765 DELB $T=654100 759480 0 0 $X=654100 $Y=759100
X1078 3766 1 2 3762 DELB $T=657820 860280 1 0 $X=657820 $Y=854860
X1079 3810 1 2 3827 DELB $T=662160 890520 0 0 $X=662160 $Y=890140
X1080 3831 1 2 3856 DELB $T=668360 799800 1 0 $X=668360 $Y=794380
X1081 3854 1 2 3869 DELB $T=672700 759480 1 0 $X=672700 $Y=754060
X1082 3917 1 2 3950 DELB $T=685100 819960 0 0 $X=685100 $Y=819580
X1083 3876 1 2 3923 DELB $T=685100 840120 1 0 $X=685100 $Y=834700
X1084 3885 1 2 3924 DELB $T=686340 729240 1 0 $X=686340 $Y=723820
X1085 3952 1 2 3980 DELB $T=690680 759480 1 0 $X=690680 $Y=754060
X1086 3905 1 2 3879 DELB $T=693160 850200 0 0 $X=693160 $Y=849820
X1087 3985 1 2 4026 DELB $T=696260 880440 0 0 $X=696260 $Y=880060
X1088 3963 1 2 3975 DELB $T=698740 729240 0 0 $X=698740 $Y=728860
X1089 3953 1 2 3976 DELB $T=699360 819960 0 0 $X=699360 $Y=819580
X1090 4015 1 2 4036 DELB $T=703700 759480 0 0 $X=703700 $Y=759100
X1091 729 1 2 4038 DELB $T=704320 729240 0 0 $X=704320 $Y=728860
X1092 3987 1 2 4043 DELB $T=704940 819960 0 0 $X=704940 $Y=819580
X1093 4008 1 2 3997 DELB $T=706180 890520 0 0 $X=706180 $Y=890140
X1094 4023 1 2 4094 DELB $T=709900 759480 1 0 $X=709900 $Y=754060
X1095 740 1 2 747 DELB $T=711140 729240 1 0 $X=711140 $Y=723820
X1096 4121 1 2 4142 DELB $T=716720 729240 1 0 $X=716720 $Y=723820
X1097 4037 1 2 4083 DELB $T=716720 779640 1 0 $X=716720 $Y=774220
X1098 4124 1 2 4131 DELB $T=718580 880440 0 0 $X=718580 $Y=880060
X1099 4113 1 2 4119 DELB $T=720440 729240 0 0 $X=720440 $Y=728860
X1100 4095 1 2 4126 DELB $T=721680 769560 0 0 $X=721680 $Y=769180
X1101 4089 1 2 4017 DELB $T=723540 840120 1 0 $X=723540 $Y=834700
X1102 763 1 2 773 DELB $T=724160 890520 0 0 $X=724160 $Y=890140
X1103 4187 1 2 4215 DELB $T=732220 890520 0 0 $X=732220 $Y=890140
X1104 785 1 2 797 DELB $T=734700 789720 1 0 $X=734700 $Y=784300
X1105 4122 1 2 4145 DELB $T=735940 749400 0 0 $X=735940 $Y=749020
X1106 4206 1 2 4210 DELB $T=735940 840120 0 0 $X=735940 $Y=839740
X1107 4076 1 2 4109 DELB $T=736560 850200 1 0 $X=736560 $Y=844780
X1108 4058 1 2 4067 DELB $T=741520 759480 1 0 $X=741520 $Y=754060
X1109 4223 1 2 4265 DELB $T=745860 809880 0 0 $X=745860 $Y=809500
X1110 4228 1 2 4273 DELB $T=747720 850200 1 0 $X=747720 $Y=844780
X1111 4231 1 2 4260 DELB $T=748340 870360 1 0 $X=748340 $Y=864940
X1112 829 1 2 4331 DELB $T=754540 749400 0 0 $X=754540 $Y=749020
X1113 4117 1 2 4141 DELB $T=755780 809880 0 0 $X=755780 $Y=809500
X1114 4373 1 2 4406 DELB $T=768180 860280 1 0 $X=768180 $Y=854860
X1115 869 1 2 879 DELB $T=775620 739320 0 0 $X=775620 $Y=738940
X1116 4443 1 2 4436 DELB $T=776860 799800 0 0 $X=776860 $Y=799420
X1117 4447 1 2 4449 DELB $T=778100 779640 1 0 $X=778100 $Y=774220
X1118 4453 1 2 4481 DELB $T=779960 870360 1 0 $X=779960 $Y=864940
X1119 880 1 2 890 DELB $T=781820 830040 1 0 $X=781820 $Y=824620
X1120 4488 1 2 4479 DELB $T=786780 870360 1 0 $X=786780 $Y=864940
X1121 4468 1 2 4541 DELB $T=789880 840120 1 0 $X=789880 $Y=834700
X1122 4513 1 2 4508 DELB $T=791120 799800 0 0 $X=791120 $Y=799420
X1123 4486 1 2 4570 DELB $T=798560 729240 0 0 $X=798560 $Y=728860
X1124 4588 1 2 4607 DELB $T=801660 739320 1 0 $X=801660 $Y=733900
X1125 4611 1 2 4644 DELB $T=805380 840120 1 0 $X=805380 $Y=834700
X1126 4629 1 2 4654 DELB $T=807860 799800 0 0 $X=807860 $Y=799420
X1127 4617 1 2 4651 DELB $T=814680 799800 0 0 $X=814680 $Y=799420
X1128 4670 1 2 4694 DELB $T=814680 840120 1 0 $X=814680 $Y=834700
X1129 4671 1 2 4695 DELB $T=814680 870360 1 0 $X=814680 $Y=864940
X1130 4643 1 2 4669 DELB $T=816540 769560 1 0 $X=816540 $Y=764140
X1131 4714 1 2 4722 DELB $T=822740 799800 0 0 $X=822740 $Y=799420
X1132 4711 1 2 4750 DELB $T=828320 759480 0 0 $X=828320 $Y=759100
X1133 4757 1 2 4787 DELB $T=829560 850200 0 0 $X=829560 $Y=849820
X1134 4779 1 2 4770 DELB $T=832660 769560 1 0 $X=832660 $Y=764140
X1135 4836 1 2 4853 DELB $T=846300 799800 0 0 $X=846300 $Y=799420
X1136 4858 1 2 4881 DELB $T=848160 860280 0 0 $X=848160 $Y=859900
X1137 4842 1 2 4845 DELB $T=853740 799800 0 0 $X=853740 $Y=799420
X1138 4907 1 2 4941 DELB $T=859940 850200 0 0 $X=859940 $Y=849820
X1139 981 1 2 986 DELB $T=861800 890520 0 0 $X=861800 $Y=890140
X1140 988 1 2 4984 DELB $T=867380 890520 0 0 $X=867380 $Y=890140
X1141 4959 1 2 993 DELB $T=868000 729240 1 0 $X=868000 $Y=723820
X1142 4994 1 2 4990 DELB $T=873580 749400 1 0 $X=873580 $Y=743980
X1143 5000 1 2 4992 DELB $T=874200 860280 1 0 $X=874200 $Y=854860
X1144 5004 1 2 5002 DELB $T=876680 759480 0 0 $X=876680 $Y=759100
X1145 5006 1 2 5035 DELB $T=876680 799800 1 0 $X=876680 $Y=794380
X1146 4993 1 2 5028 DELB $T=879780 860280 1 0 $X=879780 $Y=854860
X1147 5048 1 2 5075 DELB $T=882260 890520 0 0 $X=882260 $Y=890140
X1148 5120 1 2 5092 DELB $T=897760 819960 1 0 $X=897760 $Y=814540
X1149 5134 1 2 5164 DELB $T=898380 789720 1 0 $X=898380 $Y=784300
X1150 5115 1 2 5124 DELB $T=900240 789720 0 0 $X=900240 $Y=789340
X1151 1034 1 2 1037 DELB $T=905820 900600 1 0 $X=905820 $Y=895180
X1152 5160 1 2 5168 DELB $T=910160 739320 1 0 $X=910160 $Y=733900
X1153 5202 1 2 5209 DELB $T=911400 799800 0 0 $X=911400 $Y=799420
X1154 5216 1 2 5232 DELB $T=913880 840120 0 0 $X=913880 $Y=839740
X1155 5083 1 2 5105 DELB $T=915120 860280 0 0 $X=915120 $Y=859900
X1156 5116 1 2 5208 DELB $T=919460 779640 0 0 $X=919460 $Y=779260
X1157 5142 1 2 5188 DELB $T=919460 890520 1 0 $X=919460 $Y=885100
X1158 5165 1 2 5125 DELB $T=922560 809880 1 0 $X=922560 $Y=804460
X1159 5275 1 2 5276 DELB $T=927520 779640 0 0 $X=927520 $Y=779260
X1160 5283 1 2 5282 DELB $T=928140 809880 1 0 $X=928140 $Y=804460
X1161 5270 1 2 5277 DELB $T=931860 870360 1 0 $X=931860 $Y=864940
X1162 5268 1 2 5279 DELB $T=933100 729240 0 0 $X=933100 $Y=728860
X1163 5321 1 2 5346 DELB $T=933720 809880 1 0 $X=933720 $Y=804460
X1164 5342 1 2 5341 DELB $T=937440 759480 0 0 $X=937440 $Y=759100
X1165 1069 1 2 5419 DELB $T=943640 729240 1 0 $X=943640 $Y=723820
X1166 5410 1 2 5436 DELB $T=947360 840120 0 0 $X=947360 $Y=839740
X1167 5372 1 2 5353 DELB $T=947980 799800 0 0 $X=947980 $Y=799420
X1168 5400 1 2 5390 DELB $T=951080 870360 1 0 $X=951080 $Y=864940
X1169 5386 1 2 5426 DELB $T=952320 739320 1 0 $X=952320 $Y=733900
X1170 5465 1 2 5491 DELB $T=956040 850200 1 0 $X=956040 $Y=844780
X1171 1081 1 2 1087 DELB $T=956660 729240 1 0 $X=956660 $Y=723820
X1172 5440 1 2 5471 DELB $T=957280 830040 0 0 $X=957280 $Y=829660
X1173 5481 1 2 5387 DELB $T=958520 799800 0 0 $X=958520 $Y=799420
X1174 5479 1 2 5455 DELB $T=961620 870360 0 0 $X=961620 $Y=869980
X1175 5518 1 2 5553 DELB $T=967200 759480 0 0 $X=967200 $Y=759100
X1176 5542 1 2 5544 DELB $T=970300 809880 0 0 $X=970300 $Y=809500
X1177 5524 1 2 5545 DELB $T=974640 819960 0 0 $X=974640 $Y=819580
X1178 5534 1 2 5539 DELB $T=975260 729240 1 0 $X=975260 $Y=723820
X1179 5550 1 2 5552 DELB $T=978980 759480 1 0 $X=978980 $Y=754060
X1180 5525 1 2 5555 DELB $T=979600 830040 0 0 $X=979600 $Y=829660
X1181 5598 1 2 5626 DELB $T=982700 779640 1 0 $X=982700 $Y=774220
X1182 5612 1 2 5620 DELB $T=985800 739320 1 0 $X=985800 $Y=733900
X1183 5607 1 2 5617 DELB $T=987040 840120 1 0 $X=987040 $Y=834700
X1184 5136 1 2 5156 DELB $T=988280 870360 0 0 $X=988280 $Y=869980
X1185 5656 1 2 5672 DELB $T=992620 739320 1 0 $X=992620 $Y=733900
X1186 5660 1 2 5684 DELB $T=998820 890520 1 0 $X=998820 $Y=885100
X1187 5679 1 2 5707 DELB $T=1001300 830040 0 0 $X=1001300 $Y=829660
X1188 5744 1 2 5772 DELB $T=1009980 809880 0 0 $X=1009980 $Y=809500
X1189 5737 1 2 5773 DELB $T=1009980 830040 0 0 $X=1009980 $Y=829660
X1190 5777 1 2 5770 DELB $T=1011220 729240 0 0 $X=1011220 $Y=728860
X1191 5768 1 2 5776 DELB $T=1011840 769560 1 0 $X=1011840 $Y=764140
X1192 5812 1 2 5815 DELB $T=1018040 769560 1 0 $X=1018040 $Y=764140
X1193 5821 1 2 5858 DELB $T=1025480 840120 1 0 $X=1025480 $Y=834700
X1194 5846 1 2 5816 DELB $T=1026720 739320 0 0 $X=1026720 $Y=738940
X1195 5662 1 2 5728 DELB $T=1028580 870360 0 0 $X=1028580 $Y=869980
X1196 5907 1 2 5908 DELB $T=1033540 779640 1 0 $X=1033540 $Y=774220
X1197 5944 1 2 5915 DELB $T=1043460 739320 1 0 $X=1043460 $Y=733900
X1198 5933 1 2 5934 DELB $T=1044080 779640 1 0 $X=1044080 $Y=774220
X1199 5960 1 2 5992 DELB $T=1045940 809880 1 0 $X=1045940 $Y=804460
X1200 5990 1 2 6014 DELB $T=1049040 809880 0 0 $X=1049040 $Y=809500
X1201 5986 1 2 6022 DELB $T=1054620 749400 1 0 $X=1054620 $Y=743980
X1202 6011 1 2 6052 DELB $T=1056480 809880 1 0 $X=1056480 $Y=804460
X1203 6037 1 2 6061 DELB $T=1057720 830040 1 0 $X=1057720 $Y=824620
X1204 6016 1 2 6025 DELB $T=1058340 880440 1 0 $X=1058340 $Y=875020
X1205 6062 1 2 6070 DELB $T=1062060 850200 0 0 $X=1062060 $Y=849820
X1206 6032 1 2 6063 DELB $T=1062680 749400 1 0 $X=1062680 $Y=743980
X1207 6085 1 2 6113 DELB $T=1067020 830040 1 0 $X=1067020 $Y=824620
X1208 6075 1 2 6089 DELB $T=1067640 789720 1 0 $X=1067640 $Y=784300
X1209 6055 1 2 6096 DELB $T=1067640 880440 1 0 $X=1067640 $Y=875020
X1210 6006 1 2 5999 DELB $T=1068880 759480 1 0 $X=1068880 $Y=754060
X1211 6094 1 2 6086 DELB $T=1071360 870360 0 0 $X=1071360 $Y=869980
X1212 6172 1 2 6192 DELB $T=1084380 840120 0 0 $X=1084380 $Y=839740
X1213 1223 1 2 6177 DELB $T=1085620 729240 1 0 $X=1085620 $Y=723820
X1214 6092 1 2 6134 DELB $T=1086240 769560 1 0 $X=1086240 $Y=764140
X1215 6185 1 2 6189 DELB $T=1086860 870360 0 0 $X=1086860 $Y=869980
X1216 6165 1 2 6155 DELB $T=1089960 830040 0 0 $X=1089960 $Y=829660
X1217 6228 1 2 6258 DELB $T=1099260 789720 0 0 $X=1099260 $Y=789340
X1218 6193 1 2 6229 DELB $T=1102360 880440 1 0 $X=1102360 $Y=875020
X1219 6225 1 2 6301 DELB $T=1102980 739320 1 0 $X=1102980 $Y=733900
X1220 6227 1 2 6265 DELB $T=1106080 749400 0 0 $X=1106080 $Y=749020
X1221 6259 1 2 6292 DELB $T=1106700 729240 1 0 $X=1106700 $Y=723820
X1222 6317 1 2 6325 DELB $T=1111040 769560 1 0 $X=1111040 $Y=764140
X1223 6323 1 2 6351 DELB $T=1111040 880440 0 0 $X=1111040 $Y=880060
X1224 6302 1 2 6308 DELB $T=1124060 789720 0 0 $X=1124060 $Y=789340
X1225 1652 1 2 1653 DELA $T=277760 840120 0 0 $X=277760 $Y=839740
X1226 1881 1 2 1901 DELA $T=317440 739320 0 0 $X=317440 $Y=738940
X1227 1929 1 2 1941 DELA $T=339760 799800 1 0 $X=339760 $Y=794380
X1228 2002 1 2 2022 DELA $T=341000 809880 0 0 $X=341000 $Y=809500
X1229 2061 1 2 2095 DELA $T=345960 870360 1 0 $X=345960 $Y=864940
X1230 2100 1 2 2134 DELA $T=350920 860280 0 0 $X=350920 $Y=859900
X1231 2171 1 2 2190 DELA $T=361460 870360 1 0 $X=361460 $Y=864940
X1232 2191 1 2 2219 DELA $T=365800 870360 0 0 $X=365800 $Y=869980
X1233 2206 1 2 2235 DELA $T=368280 819960 1 0 $X=368280 $Y=814540
X1234 2200 1 2 2244 DELA $T=375720 830040 1 0 $X=375720 $Y=824620
X1235 251 1 2 256 DELA $T=380060 900600 1 0 $X=380060 $Y=895180
X1236 2287 1 2 2318 DELA $T=380680 830040 1 0 $X=380680 $Y=824620
X1237 2321 1 2 2352 DELA $T=385020 900600 1 0 $X=385020 $Y=895180
X1238 2349 1 2 2377 DELA $T=388740 819960 0 0 $X=388740 $Y=819580
X1239 2383 1 2 2408 DELA $T=394320 809880 1 0 $X=394320 $Y=804460
X1240 2411 1 2 2439 DELA $T=399280 799800 1 0 $X=399280 $Y=794380
X1241 284 1 2 289 DELA $T=404240 799800 1 0 $X=404240 $Y=794380
X1242 2442 1 2 2478 DELA $T=404860 890520 1 0 $X=404860 $Y=885100
X1243 2483 1 2 2509 DELA $T=409820 890520 1 0 $X=409820 $Y=885100
X1244 2550 1 2 2573 DELA $T=422220 870360 1 0 $X=422220 $Y=864940
X1245 2561 1 2 2581 DELA $T=424700 769560 0 0 $X=424700 $Y=769180
X1246 2586 1 2 2608 DELA $T=429660 860280 0 0 $X=429660 $Y=859900
X1247 319 1 2 326 DELA $T=431520 769560 1 0 $X=431520 $Y=764140
X1248 2597 1 2 2617 DELA $T=432140 789720 1 0 $X=432140 $Y=784300
X1249 2615 1 2 2640 DELA $T=436480 769560 1 0 $X=436480 $Y=764140
X1250 2662 1 2 2698 DELA $T=445160 759480 0 0 $X=445160 $Y=759100
X1251 2718 1 2 2737 DELA $T=453840 739320 1 0 $X=453840 $Y=733900
X1252 408 1 2 416 DELA $T=500340 890520 1 0 $X=500340 $Y=885100
X1253 2924 1 2 2948 DELA $T=501580 850200 1 0 $X=501580 $Y=844780
X1254 2989 1 2 3014 DELA $T=505920 739320 1 0 $X=505920 $Y=733900
X1255 3019 1 2 3039 DELA $T=510880 739320 1 0 $X=510880 $Y=733900
X1256 3029 1 2 3005 DELA $T=512740 850200 1 0 $X=512740 $Y=844780
X1257 3184 1 2 3255 DELA $T=556140 729240 0 0 $X=556140 $Y=728860
X1258 3284 1 2 3310 DELA $T=561720 729240 0 0 $X=561720 $Y=728860
X1259 489 1 2 496 DELA $T=567300 729240 1 0 $X=567300 $Y=723820
X1260 3342 1 2 3366 DELA $T=571640 729240 0 0 $X=571640 $Y=728860
X1261 518 1 2 530 DELA $T=583420 729240 1 0 $X=583420 $Y=723820
X1262 3346 1 2 3277 DELA $T=584660 809880 1 0 $X=584660 $Y=804460
X1263 3438 1 2 3439 DELA $T=590240 759480 1 0 $X=590240 $Y=754060
X1264 3502 1 2 3542 DELA $T=608220 789720 1 0 $X=608220 $Y=784300
X1265 3547 1 2 3565 DELA $T=610080 749400 0 0 $X=610080 $Y=749020
X1266 3588 1 2 3615 DELA $T=618140 840120 0 0 $X=618140 $Y=839740
X1267 3586 1 2 3570 DELA $T=628060 779640 1 0 $X=628060 $Y=774220
X1268 3703 1 2 3725 DELA $T=641700 860280 1 0 $X=641700 $Y=854860
X1269 4227 1 2 4238 DELA $T=740900 809880 0 0 $X=740900 $Y=809500
X1270 4217 1 2 4237 DELA $T=750820 809880 0 0 $X=750820 $Y=809500
X1271 4416 1 2 4457 DELA $T=780580 739320 0 0 $X=780580 $Y=738940
X1272 4511 1 2 4543 DELA $T=793600 769560 1 0 $X=793600 $Y=764140
X1273 4536 1 2 4550 DELA $T=795460 870360 0 0 $X=795460 $Y=869980
X1274 4749 1 2 4781 DELA $T=828940 880440 1 0 $X=828940 $Y=875020
X1275 5444 1 2 5478 DELA $T=953560 799800 0 0 $X=953560 $Y=799420
X1276 5469 1 2 5500 DELA $T=983320 809880 0 0 $X=983320 $Y=809500
X1277 5790 1 2 5791 DELA $T=1013700 870360 0 0 $X=1013700 $Y=869980
X1278 5806 1 2 5799 DELA $T=1016800 840120 1 0 $X=1016800 $Y=834700
X1279 5841 1 2 5843 DELA $T=1024240 749400 1 0 $X=1024240 $Y=743980
X1280 5847 1 2 5833 DELA $T=1024860 779640 1 0 $X=1024860 $Y=774220
X1281 5784 1 2 5785 DELA $T=1031680 789720 1 0 $X=1031680 $Y=784300
X1282 5897 1 2 5916 DELA $T=1032300 749400 1 0 $X=1032300 $Y=743980
X1283 5909 1 2 5899 DELA $T=1039120 769560 0 0 $X=1039120 $Y=769180
X1284 5929 1 2 5951 DELA $T=1040980 880440 1 0 $X=1040980 $Y=875020
X1285 1315 7 1371 2 1 1394 QDFFRBN $T=221340 749400 0 0 $X=221340 $Y=749020
X1286 1363 7 1371 2 1 19 QDFFRBN $T=228160 749400 1 0 $X=228160 $Y=743980
X1287 1441 7 1371 2 1 25 QDFFRBN $T=239320 739320 0 0 $X=239320 $Y=738940
X1288 1471 7 1371 2 1 1495 QDFFRBN $T=244900 729240 0 0 $X=244900 $Y=728860
X1289 1528 7 1487 2 1 35 QDFFRBN $T=256680 850200 1 180 $X=244900 $Y=849820
X1290 1557 7 1487 2 1 1429 QDFFRBN $T=256680 860280 0 180 $X=244900 $Y=854860
X1291 68 7 48 2 1 43 QDFFRBN $T=262260 729240 0 180 $X=250480 $Y=723820
X1292 1573 7 1487 2 1 37 QDFFRBN $T=264740 850200 0 180 $X=252960 $Y=844780
X1293 1579 7 1487 2 1 1520 QDFFRBN $T=266600 840120 0 180 $X=254820 $Y=834700
X1294 57 7 1371 2 1 70 QDFFRBN $T=259160 729240 0 0 $X=259160 $Y=728860
X1295 1577 7 1608 2 1 1635 QDFFRBN $T=262880 819960 0 0 $X=262880 $Y=819580
X1296 1578 7 1487 2 1 1452 QDFFRBN $T=262880 830040 0 0 $X=262880 $Y=829660
X1297 1604 7 1487 2 1 1453 QDFFRBN $T=275900 850200 1 180 $X=264120 $Y=849820
X1298 1588 7 75 2 1 81 QDFFRBN $T=264740 729240 1 0 $X=264740 $Y=723820
X1299 1667 7 1608 2 1 53 QDFFRBN $T=281480 850200 0 180 $X=269700 $Y=844780
X1300 1682 7 1608 2 1 72 QDFFRBN $T=282720 840120 0 180 $X=270940 $Y=834700
X1301 1717 7 1608 2 1 79 QDFFRBN $T=288300 830040 1 180 $X=276520 $Y=829660
X1302 1641 7 1714 2 1 1712 QDFFRBN $T=281480 830040 1 0 $X=281480 $Y=824620
X1303 1695 7 1608 2 1 1612 QDFFRBN $T=283340 819960 0 0 $X=283340 $Y=819580
X1304 1747 7 1714 2 1 1678 QDFFRBN $T=295120 850200 0 180 $X=283340 $Y=844780
X1305 1687 7 75 2 1 1809 QDFFRBN $T=289540 729240 0 0 $X=289540 $Y=728860
X1306 1782 7 1714 2 1 109 QDFFRBN $T=307520 840120 1 180 $X=295740 $Y=839740
X1307 1798 7 1824 2 1 1814 QDFFRBN $T=300700 809880 1 0 $X=300700 $Y=804460
X1308 1757 7 1824 2 1 1794 QDFFRBN $T=300700 819960 1 0 $X=300700 $Y=814540
X1309 1898 7 75 2 1 1847 QDFFRBN $T=321780 749400 1 180 $X=310000 $Y=749020
X1310 1931 7 138 2 1 1607 QDFFRBN $T=322400 749400 0 180 $X=310620 $Y=743980
X1311 1876 7 1873 2 1 1823 QDFFRBN $T=324260 819960 1 180 $X=312480 $Y=819580
X1312 1905 7 120 2 1 132 QDFFRBN $T=324260 850200 0 180 $X=312480 $Y=844780
X1313 1906 7 1824 2 1 1580 QDFFRBN $T=324880 809880 1 180 $X=313100 $Y=809500
X1314 1907 7 1878 2 1 134 QDFFRBN $T=324880 830040 1 180 $X=313100 $Y=829660
X1315 1925 7 1878 2 1 139 QDFFRBN $T=325500 840120 1 180 $X=313720 $Y=839740
X1316 1939 7 1824 2 1 1613 QDFFRBN $T=326120 799800 1 180 $X=314340 $Y=799420
X1317 1932 7 1873 2 1 1599 QDFFRBN $T=328600 819960 0 180 $X=316820 $Y=814540
X1318 1956 1935 1873 2 1 1882 QDFFRBN $T=329220 830040 0 180 $X=317440 $Y=824620
X1319 1946 7 120 2 1 1849 QDFFRBN $T=330460 850200 1 180 $X=318680 $Y=849820
X1320 2025 1935 1873 2 1 1564 QDFFRBN $T=341620 819960 0 180 $X=329840 $Y=814540
X1321 1985 1935 1970 2 1 1997 QDFFRBN $T=334180 830040 1 0 $X=334180 $Y=824620
X1322 2109 1935 2054 2 1 1984 QDFFRBN $T=353400 819960 0 180 $X=341620 $Y=814540
X1323 2110 1935 1970 2 1 1996 QDFFRBN $T=353400 840120 0 180 $X=341620 $Y=834700
X1324 2069 1935 2054 2 1 2073 QDFFRBN $T=346580 830040 0 0 $X=346580 $Y=829660
X1325 2174 1935 2054 2 1 2122 QDFFRBN $T=365180 819960 0 180 $X=353400 $Y=814540
X1326 2195 1935 2054 2 1 176 QDFFRBN $T=367660 840120 0 180 $X=355880 $Y=834700
X1327 2185 1935 2164 2 1 2151 QDFFRBN $T=369520 830040 0 180 $X=357740 $Y=824620
X1328 2229 1935 2182 2 1 144 QDFFRBN $T=373240 850200 0 180 $X=361460 $Y=844780
X1329 2253 1935 2182 2 1 1855 QDFFRBN $T=376340 840120 1 180 $X=364560 $Y=839740
X1330 2240 1935 2182 2 1 209 QDFFRBN $T=378200 850200 1 180 $X=366420 $Y=849820
X1331 2316 1935 2182 2 1 2227 QDFFRBN $T=383160 840120 0 180 $X=371380 $Y=834700
X1332 2309 1935 2182 2 1 217 QDFFRBN $T=385020 860280 0 180 $X=373240 $Y=854860
X1333 2327 1935 2164 2 1 2250 QDFFRBN $T=387500 819960 1 180 $X=375720 $Y=819580
X1334 2314 1935 2373 2 1 1886 QDFFRBN $T=384400 850200 0 0 $X=384400 $Y=849820
X1335 2348 258 2373 2 1 2397 QDFFRBN $T=388120 870360 1 0 $X=388120 $Y=864940
X1336 2496 258 2373 2 1 227 QDFFRBN $T=412920 870360 0 180 $X=401140 $Y=864940
X1337 2395 1935 2164 2 1 2400 QDFFRBN $T=414160 819960 0 180 $X=402380 $Y=814540
X1338 2512 258 2373 2 1 2161 QDFFRBN $T=416020 870360 1 180 $X=404240 $Y=869980
X1339 2393 1935 2514 2 1 2476 QDFFRBN $T=409820 830040 0 0 $X=409820 $Y=829660
X1340 2402 1935 2514 2 1 2506 QDFFRBN $T=411680 850200 1 0 $X=411680 $Y=844780
X1341 2567 1935 2532 2 1 1860 QDFFRBN $T=426560 809880 1 180 $X=414780 $Y=809500
X1342 2572 1935 2514 2 1 2494 QDFFRBN $T=428420 850200 1 180 $X=416640 $Y=849820
X1343 2555 258 2545 2 1 2403 QDFFRBN $T=429040 880440 0 180 $X=417260 $Y=875020
X1344 2562 1935 2514 2 1 2329 QDFFRBN $T=429660 860280 0 180 $X=417880 $Y=854860
X1345 2582 1935 2514 2 1 1893 QDFFRBN $T=432140 840120 1 180 $X=420360 $Y=839740
X1346 2591 1935 2532 2 1 2597 QDFFRBN $T=429660 809880 1 0 $X=429660 $Y=804460
X1347 2587 1935 2532 2 1 2645 QDFFRBN $T=429660 830040 1 0 $X=429660 $Y=824620
X1348 2593 1935 2620 2 1 2643 QDFFRBN $T=430280 779640 0 0 $X=430280 $Y=779260
X1349 2606 258 2545 2 1 2420 QDFFRBN $T=442060 870360 1 180 $X=430280 $Y=869980
X1350 2629 258 2545 2 1 2211 QDFFRBN $T=442680 880440 0 180 $X=430900 $Y=875020
X1351 2592 1935 2545 2 1 2223 QDFFRBN $T=443300 850200 1 180 $X=431520 $Y=849820
X1352 2600 1935 2532 2 1 2559 QDFFRBN $T=432140 819960 1 0 $X=432140 $Y=814540
X1353 2604 258 335 2 1 2676 QDFFRBN $T=432760 890520 0 0 $X=432760 $Y=890140
X1354 2611 1935 2632 2 1 2669 QDFFRBN $T=434620 840120 0 0 $X=434620 $Y=839740
X1355 2613 1935 2632 2 1 2602 QDFFRBN $T=435240 850200 1 0 $X=435240 $Y=844780
X1356 2623 1935 2632 2 1 2483 QDFFRBN $T=437100 860280 1 0 $X=437100 $Y=854860
X1357 2657 258 2710 2 1 2720 QDFFRBN $T=443300 870360 0 0 $X=443300 $Y=869980
X1358 2661 1935 2667 2 1 2704 QDFFRBN $T=443920 769560 0 0 $X=443920 $Y=769180
X1359 2664 258 2710 2 1 2552 QDFFRBN $T=444540 880440 1 0 $X=444540 $Y=875020
X1360 2730 1935 2697 2 1 2499 QDFFRBN $T=458800 819960 0 180 $X=447020 $Y=814540
X1361 2681 1935 2725 2 1 2709 QDFFRBN $T=447020 850200 0 0 $X=447020 $Y=849820
X1362 2685 258 356 2 1 2740 QDFFRBN $T=447640 880440 0 0 $X=447640 $Y=880060
X1363 343 258 335 2 1 2741 QDFFRBN $T=447640 890520 0 0 $X=447640 $Y=890140
X1364 2696 1935 2697 2 1 2724 QDFFRBN $T=448880 809880 0 0 $X=448880 $Y=809500
X1365 2707 1935 2667 2 1 2729 QDFFRBN $T=450740 779640 1 0 $X=450740 $Y=774220
X1366 2766 1935 2697 2 1 2628 QDFFRBN $T=465000 840120 0 180 $X=453220 $Y=834700
X1367 2748 1935 2632 2 1 2716 QDFFRBN $T=465000 860280 1 180 $X=453220 $Y=859900
X1368 2723 1935 2667 2 1 2759 QDFFRBN $T=454460 789720 1 0 $X=454460 $Y=784300
X1369 2726 258 356 2 1 2721 QDFFRBN $T=455080 870360 0 0 $X=455080 $Y=869980
X1370 2734 1935 2725 2 1 2804 QDFFRBN $T=456320 840120 0 0 $X=456320 $Y=839740
X1371 2738 1935 2782 2 1 2789 QDFFRBN $T=458180 769560 0 0 $X=458180 $Y=769180
X1372 2777 2796 2667 2 1 2744 QDFFRBN $T=471200 799800 1 180 $X=459420 $Y=799420
X1373 2752 1935 2797 2 1 2411 QDFFRBN $T=460660 819960 1 0 $X=460660 $Y=814540
X1374 2823 258 356 2 1 2757 QDFFRBN $T=473680 900600 0 180 $X=461900 $Y=895180
X1375 2767 1935 2797 2 1 2627 QDFFRBN $T=463140 809880 0 0 $X=463140 $Y=809500
X1376 2768 1935 2725 2 1 2827 QDFFRBN $T=463140 850200 0 0 $X=463140 $Y=849820
X1377 2772 1935 2797 2 1 2835 QDFFRBN $T=464380 819960 0 0 $X=464380 $Y=819580
X1378 2825 1935 2782 2 1 2543 QDFFRBN $T=477400 759480 1 180 $X=465620 $Y=759100
X1379 2788 1935 2710 2 1 2859 QDFFRBN $T=466860 860280 1 0 $X=466860 $Y=854860
X1380 2791 1935 2710 2 1 2847 QDFFRBN $T=467480 870360 1 0 $X=467480 $Y=864940
X1381 2803 1935 2842 2 1 2822 QDFFRBN $T=469340 759480 1 0 $X=469340 $Y=754060
X1382 2851 258 371 2 1 2746 QDFFRBN $T=481120 890520 1 180 $X=469340 $Y=890140
X1383 2809 1935 2842 2 1 2861 QDFFRBN $T=470580 749400 1 0 $X=470580 $Y=743980
X1384 2810 1935 2842 2 1 2718 QDFFRBN $T=470580 749400 0 0 $X=470580 $Y=749020
X1385 2802 1935 2725 2 1 2850 QDFFRBN $T=470580 850200 1 0 $X=470580 $Y=844780
X1386 2854 2796 2782 2 1 2806 QDFFRBN $T=483600 779640 0 180 $X=471820 $Y=774220
X1387 2865 2796 2782 2 1 2818 QDFFRBN $T=484220 769560 1 180 $X=472440 $Y=769180
X1388 2826 2796 2782 2 1 2668 QDFFRBN $T=484220 799800 1 180 $X=472440 $Y=799420
X1389 2829 2796 2797 2 1 2884 QDFFRBN $T=474300 819960 1 0 $X=474300 $Y=814540
X1390 2834 258 2828 2 1 2442 QDFFRBN $T=474920 870360 0 0 $X=474920 $Y=869980
X1391 2878 2796 2797 2 1 2840 QDFFRBN $T=488560 819960 1 180 $X=476780 $Y=819580
X1392 2844 2796 2725 2 1 2880 QDFFRBN $T=477400 850200 0 0 $X=477400 $Y=849820
X1393 2862 2796 2725 2 1 2889 QDFFRBN $T=481740 840120 0 0 $X=481740 $Y=839740
X1394 2912 2796 2828 2 1 388 QDFFRBN $T=493520 860280 0 180 $X=481740 $Y=854860
X1395 2868 393 2842 2 1 2916 QDFFRBN $T=482980 759480 1 0 $X=482980 $Y=754060
X1396 2869 2796 2797 2 1 2892 QDFFRBN $T=482980 809880 1 0 $X=482980 $Y=804460
X1397 2870 258 371 2 1 2908 QDFFRBN $T=482980 890520 0 0 $X=482980 $Y=890140
X1398 2911 393 392 2 1 2792 QDFFRBN $T=496000 739320 0 180 $X=484220 $Y=733900
X1399 2873 393 2842 2 1 2934 QDFFRBN $T=484220 759480 0 0 $X=484220 $Y=759100
X1400 395 393 392 2 1 387 QDFFRBN $T=484840 729240 1 0 $X=484840 $Y=723820
X1401 2877 2796 2902 2 1 2928 QDFFRBN $T=485460 779640 0 0 $X=485460 $Y=779260
X1402 2961 393 2902 2 1 2881 QDFFRBN $T=498480 769560 1 180 $X=486700 $Y=769180
X1403 2938 258 2907 2 1 2886 QDFFRBN $T=499100 880440 0 180 $X=487320 $Y=875020
X1404 2900 2796 2930 2 1 2924 QDFFRBN $T=488560 809880 0 0 $X=488560 $Y=809500
X1405 2946 2796 2828 2 1 2897 QDFFRBN $T=500340 870360 0 180 $X=488560 $Y=864940
X1406 2909 2796 2947 2 1 2979 QDFFRBN $T=491040 799800 1 0 $X=491040 $Y=794380
X1407 2927 2796 2966 2 1 2610 QDFFRBN $T=495380 840120 0 0 $X=495380 $Y=839740
X1408 2935 393 2986 2 1 421 QDFFRBN $T=497240 729240 0 0 $X=497240 $Y=728860
X1409 2932 258 2907 2 1 3001 QDFFRBN $T=497240 890520 0 0 $X=497240 $Y=890140
X1410 2942 2796 2947 2 1 2920 QDFFRBN $T=499100 830040 1 0 $X=499100 $Y=824620
X1411 2955 2796 2966 2 1 2355 QDFFRBN $T=510880 850200 1 180 $X=499100 $Y=849820
X1412 2958 393 3010 2 1 2981 QDFFRBN $T=500960 769560 0 0 $X=500960 $Y=769180
X1413 2962 2796 2966 2 1 2988 QDFFRBN $T=500960 819960 1 0 $X=500960 $Y=814540
X1414 2975 2796 2966 2 1 2944 QDFFRBN $T=504680 860280 1 0 $X=504680 $Y=854860
X1415 2995 258 3034 2 1 3031 QDFFRBN $T=505920 870360 0 0 $X=505920 $Y=869980
X1416 3002 2796 3010 2 1 3056 QDFFRBN $T=507780 779640 0 0 $X=507780 $Y=779260
X1417 3012 393 2986 2 1 3071 QDFFRBN $T=509640 749400 0 0 $X=509640 $Y=749020
X1418 3063 2796 2966 2 1 2251 QDFFRBN $T=521420 840120 1 180 $X=509640 $Y=839740
X1419 3016 2796 2947 2 1 3048 QDFFRBN $T=510260 809880 1 0 $X=510260 $Y=804460
X1420 3020 2796 2947 2 1 3029 QDFFRBN $T=510880 830040 1 0 $X=510880 $Y=824620
X1421 3024 393 3060 2 1 3042 QDFFRBN $T=511500 729240 0 0 $X=511500 $Y=728860
X1422 3025 393 3060 2 1 3076 QDFFRBN $T=511500 739320 0 0 $X=511500 $Y=738940
X1423 3082 2796 3041 2 1 2992 QDFFRBN $T=524520 830040 1 180 $X=512740 $Y=829660
X1424 3040 258 431 2 1 3013 QDFFRBN $T=525140 890520 1 180 $X=513360 $Y=890140
X1425 432 393 3060 2 1 438 QDFFRBN $T=515840 729240 1 0 $X=515840 $Y=723820
X1426 3046 258 431 2 1 2550 QDFFRBN $T=527620 890520 0 180 $X=515840 $Y=885100
X1427 3047 2796 3010 2 1 3059 QDFFRBN $T=517080 769560 0 0 $X=517080 $Y=769180
X1428 3107 258 3034 2 1 3051 QDFFRBN $T=529480 870360 1 180 $X=517700 $Y=869980
X1429 3119 2796 3010 2 1 3065 QDFFRBN $T=531960 779640 0 180 $X=520180 $Y=774220
X1430 3079 2796 2902 2 1 3114 QDFFRBN $T=522040 809880 0 0 $X=522040 $Y=809500
X1431 3081 2796 3041 2 1 3105 QDFFRBN $T=522660 819960 1 0 $X=522660 $Y=814540
X1432 3083 2796 3034 2 1 2398 QDFFRBN $T=522660 870360 1 0 $X=522660 $Y=864940
X1433 3089 393 3135 2 1 3154 QDFFRBN $T=523900 769560 1 0 $X=523900 $Y=764140
X1434 3163 393 3118 2 1 3075 QDFFRBN $T=537540 739320 0 180 $X=525760 $Y=733900
X1435 3103 2796 3041 2 1 3147 QDFFRBN $T=525760 840120 1 0 $X=525760 $Y=834700
X1436 3150 258 431 2 1 3121 QDFFRBN $T=540640 890520 0 180 $X=528860 $Y=885100
X1437 3164 2796 3157 2 1 2383 QDFFRBN $T=543740 799800 0 180 $X=531960 $Y=794380
X1438 3143 2796 3135 2 1 3176 QDFFRBN $T=532580 769560 0 0 $X=532580 $Y=769180
X1439 3172 2796 3157 2 1 2989 QDFFRBN $T=545600 809880 1 180 $X=533820 $Y=809500
X1440 3158 457 431 2 1 441 QDFFRBN $T=546220 900600 0 180 $X=534440 $Y=895180
X1441 3175 2796 3157 2 1 3122 QDFFRBN $T=546840 819960 1 180 $X=535060 $Y=819580
X1442 3194 2796 3034 2 1 3132 QDFFRBN $T=546840 860280 1 180 $X=535060 $Y=859900
X1443 3171 2796 3135 2 1 3145 QDFFRBN $T=547460 779640 1 180 $X=535680 $Y=779260
X1444 3166 2796 3034 2 1 3078 QDFFRBN $T=547460 870360 1 180 $X=535680 $Y=869980
X1445 3200 393 3135 2 1 3170 QDFFRBN $T=549320 769560 0 180 $X=537540 $Y=764140
X1446 3179 393 3118 2 1 453 QDFFRBN $T=539400 739320 1 0 $X=539400 $Y=733900
X1447 3201 2796 3141 2 1 3139 QDFFRBN $T=551180 850200 0 180 $X=539400 $Y=844780
X1448 3188 2796 3196 2 1 3129 QDFFRBN $T=551800 830040 0 180 $X=540020 $Y=824620
X1449 3221 2796 3199 2 1 3088 QDFFRBN $T=552420 789720 1 180 $X=540640 $Y=789340
X1450 3191 457 3141 2 1 3242 QDFFRBN $T=541880 880440 0 0 $X=541880 $Y=880060
X1451 456 393 444 2 1 468 QDFFRBN $T=542500 729240 1 0 $X=542500 $Y=723820
X1452 3195 457 3141 2 1 470 QDFFRBN $T=542500 880440 1 0 $X=542500 $Y=875020
X1453 3198 2796 3223 2 1 3219 QDFFRBN $T=543120 779640 1 0 $X=543120 $Y=774220
X1454 3212 2796 3227 2 1 3249 QDFFRBN $T=548080 860280 1 0 $X=548080 $Y=854860
X1455 3216 2796 3227 2 1 3209 QDFFRBN $T=548700 860280 0 0 $X=548700 $Y=859900
X1456 3260 2796 3157 2 1 3222 QDFFRBN $T=561720 809880 1 180 $X=549940 $Y=809500
X1457 3230 393 3223 2 1 3276 QDFFRBN $T=550560 769560 1 0 $X=550560 $Y=764140
X1458 3232 2796 3227 2 1 3289 QDFFRBN $T=551180 850200 0 0 $X=551180 $Y=849820
X1459 3236 393 3118 2 1 3273 QDFFRBN $T=552420 739320 0 0 $X=552420 $Y=738940
X1460 3237 393 3118 2 1 3279 QDFFRBN $T=552420 749400 1 0 $X=552420 $Y=743980
X1461 3238 2796 3227 2 1 3278 QDFFRBN $T=552420 850200 1 0 $X=552420 $Y=844780
X1462 3241 2796 3196 2 1 3266 QDFFRBN $T=553040 830040 1 0 $X=553040 $Y=824620
X1463 3251 457 3291 2 1 2493 QDFFRBN $T=554280 880440 1 0 $X=554280 $Y=875020
X1464 3239 393 3223 2 1 462 QDFFRBN $T=567300 759480 0 180 $X=555520 $Y=754060
X1465 3261 2796 3223 2 1 3206 QDFFRBN $T=559240 789720 1 0 $X=559240 $Y=784300
X1466 3327 3314 3283 2 1 3269 QDFFRBN $T=571020 799800 1 180 $X=559240 $Y=799420
X1467 3338 3314 3223 2 1 3292 QDFFRBN $T=574740 779640 0 180 $X=562960 $Y=774220
X1468 3303 2796 3196 2 1 3346 QDFFRBN $T=563580 819960 0 0 $X=563580 $Y=819580
X1469 3305 457 3350 2 1 3218 QDFFRBN $T=564200 890520 1 0 $X=564200 $Y=885100
X1470 3306 3314 3135 2 1 504 QDFFRBN $T=564820 769560 0 0 $X=564820 $Y=769180
X1471 3367 393 490 2 1 3019 QDFFRBN $T=577840 739320 1 180 $X=566060 $Y=738940
X1472 3311 393 490 2 1 3355 QDFFRBN $T=566060 749400 1 0 $X=566060 $Y=743980
X1473 3359 3314 3283 2 1 3312 QDFFRBN $T=577840 809880 1 180 $X=566060 $Y=809500
X1474 3308 2796 3196 2 1 3336 QDFFRBN $T=566060 830040 1 0 $X=566060 $Y=824620
X1475 3371 457 3291 2 1 3313 QDFFRBN $T=577840 880440 0 180 $X=566060 $Y=875020
X1476 3388 393 490 2 1 491 QDFFRBN $T=580320 739320 0 180 $X=568540 $Y=733900
X1477 3349 3314 3397 2 1 2727 QDFFRBN $T=571640 850200 0 0 $X=571640 $Y=849820
X1478 501 457 3350 2 1 522 QDFFRBN $T=572880 900600 1 0 $X=572880 $Y=895180
X1479 3354 457 3350 2 1 3409 QDFFRBN $T=573500 890520 0 0 $X=573500 $Y=890140
X1480 3376 3314 3385 2 1 3353 QDFFRBN $T=577840 850200 1 0 $X=577840 $Y=844780
X1481 3390 3314 3385 2 1 3398 QDFFRBN $T=578460 840120 0 0 $X=578460 $Y=839740
X1482 3443 3314 3283 2 1 3399 QDFFRBN $T=591480 809880 1 180 $X=579700 $Y=809500
X1483 3437 3314 3385 2 1 3402 QDFFRBN $T=591480 830040 0 180 $X=579700 $Y=824620
X1484 3405 3314 3385 2 1 515 QDFFRBN $T=592100 819960 1 180 $X=580320 $Y=819580
X1485 3411 393 3418 2 1 3381 QDFFRBN $T=580940 749400 0 0 $X=580940 $Y=749020
X1486 3451 3314 3419 2 1 508 QDFFRBN $T=593960 779640 1 180 $X=582180 $Y=779260
X1487 3421 3314 3350 2 1 2321 QDFFRBN $T=595820 880440 0 180 $X=584040 $Y=875020
X1488 3466 3314 3418 2 1 3392 QDFFRBN $T=597060 759480 1 180 $X=585280 $Y=759100
X1489 3444 3314 3419 2 1 2615 QDFFRBN $T=598300 799800 0 180 $X=586520 $Y=794380
X1490 3476 3314 3397 2 1 2586 QDFFRBN $T=598300 870360 1 180 $X=586520 $Y=869980
X1491 3478 393 3418 2 1 499 QDFFRBN $T=598920 739320 1 180 $X=587140 $Y=738940
X1492 3479 3314 3397 2 1 3433 QDFFRBN $T=598920 860280 0 180 $X=587140 $Y=854860
X1493 3503 457 3350 2 1 2533 QDFFRBN $T=598920 890520 0 180 $X=587140 $Y=885100
X1494 3425 393 3418 2 1 523 QDFFRBN $T=600160 729240 0 180 $X=588380 $Y=723820
X1495 3435 393 3418 2 1 528 QDFFRBN $T=600780 739320 0 180 $X=589000 $Y=733900
X1496 3483 3314 3458 2 1 3449 QDFFRBN $T=603880 809880 1 180 $X=592100 $Y=809500
X1497 3516 3314 3419 2 1 526 QDFFRBN $T=604500 779640 0 180 $X=592720 $Y=774220
X1498 3518 3314 3419 2 1 3375 QDFFRBN $T=605120 769560 1 180 $X=593340 $Y=769180
X1499 3488 3314 3458 2 1 3455 QDFFRBN $T=605120 830040 0 180 $X=593340 $Y=824620
X1500 3470 393 3519 2 1 3513 QDFFRBN $T=595820 749400 1 0 $X=595820 $Y=743980
X1501 3540 3314 3510 2 1 3489 QDFFRBN $T=610700 850200 1 180 $X=598920 $Y=849820
X1502 3496 3314 3430 2 1 558 QDFFRBN $T=600160 759480 0 0 $X=600160 $Y=759100
X1503 548 550 3544 2 1 561 QDFFRBN $T=601400 729240 1 0 $X=601400 $Y=723820
X1504 3506 3314 3458 2 1 3500 QDFFRBN $T=601400 809880 1 0 $X=601400 $Y=804460
X1505 3515 550 3544 2 1 3564 QDFFRBN $T=602640 739320 1 0 $X=602640 $Y=733900
X1506 3548 3314 3510 2 1 3456 QDFFRBN $T=614420 870360 1 180 $X=602640 $Y=869980
X1507 3508 3314 3430 2 1 2751 QDFFRBN $T=603880 799800 1 0 $X=603880 $Y=794380
X1508 3522 3314 3555 2 1 3569 QDFFRBN $T=603880 809880 0 0 $X=603880 $Y=809500
X1509 3561 3314 3510 2 1 3521 QDFFRBN $T=615660 870360 0 180 $X=603880 $Y=864940
X1510 3526 3314 3430 2 1 566 QDFFRBN $T=604500 769560 1 0 $X=604500 $Y=764140
X1511 3531 457 562 2 1 3525 QDFFRBN $T=605120 890520 0 0 $X=605120 $Y=890140
X1512 3524 3314 3458 2 1 3492 QDFFRBN $T=618140 840120 0 180 $X=606360 $Y=834700
X1513 3512 457 562 2 1 552 QDFFRBN $T=606360 900600 1 0 $X=606360 $Y=895180
X1514 3537 3314 3430 2 1 3586 QDFFRBN $T=606980 769560 0 0 $X=606980 $Y=769180
X1515 3538 3314 3430 2 1 574 QDFFRBN $T=606980 779640 0 0 $X=606980 $Y=779260
X1516 3514 3314 3458 2 1 3497 QDFFRBN $T=618760 819960 1 180 $X=606980 $Y=819580
X1517 3535 3314 3385 2 1 3342 QDFFRBN $T=618760 830040 0 180 $X=606980 $Y=824620
X1518 3541 550 3519 2 1 3568 QDFFRBN $T=608220 749400 1 0 $X=608220 $Y=743980
X1519 3550 3314 3555 2 1 3559 QDFFRBN $T=610700 799800 0 0 $X=610700 $Y=799420
X1520 3605 3314 3510 2 1 2601 QDFFRBN $T=623720 850200 0 180 $X=611940 $Y=844780
X1521 3556 3314 3592 2 1 549 QDFFRBN $T=611940 850200 0 0 $X=611940 $Y=849820
X1522 3558 3314 3458 2 1 3502 QDFFRBN $T=624960 830040 1 180 $X=613180 $Y=829660
X1523 3626 3314 3510 2 1 3517 QDFFRBN $T=626820 860280 1 180 $X=615040 $Y=859900
X1524 3576 550 3519 2 1 3547 QDFFRBN $T=616280 739320 1 0 $X=616280 $Y=733900
X1525 3616 3314 3592 2 1 3423 QDFFRBN $T=628060 870360 1 180 $X=616280 $Y=869980
X1526 3648 3314 3592 2 1 535 QDFFRBN $T=630540 860280 0 180 $X=618760 $Y=854860
X1527 3587 3314 3592 2 1 3574 QDFFRBN $T=619380 819960 0 0 $X=619380 $Y=819580
X1528 3557 457 577 2 1 2561 QDFFRBN $T=631780 890520 0 180 $X=620000 $Y=885100
X1529 3598 550 3641 2 1 584 QDFFRBN $T=620620 749400 1 0 $X=620620 $Y=743980
X1530 3614 3314 3654 2 1 595 QDFFRBN $T=622480 830040 1 0 $X=622480 $Y=824620
X1531 3622 3314 3657 2 1 602 QDFFRBN $T=623100 840120 0 0 $X=623100 $Y=839740
X1532 3668 3314 3555 2 1 3624 QDFFRBN $T=635500 809880 0 180 $X=623720 $Y=804460
X1533 3578 457 577 2 1 2549 QDFFRBN $T=636120 880440 1 180 $X=624340 $Y=880060
X1534 3649 550 3644 2 1 585 QDFFRBN $T=637360 769560 1 180 $X=625580 $Y=769180
X1535 586 457 3667 2 1 611 QDFFRBN $T=625580 900600 1 0 $X=625580 $Y=895180
X1536 3663 3314 3644 2 1 3602 QDFFRBN $T=637980 779640 1 180 $X=626200 $Y=779260
X1537 3659 3314 3644 2 1 581 QDFFRBN $T=640460 789720 1 180 $X=628680 $Y=789340
X1538 3685 550 3641 2 1 3634 QDFFRBN $T=641080 759480 0 180 $X=629300 $Y=754060
X1539 3681 550 3519 2 1 3610 QDFFRBN $T=641700 739320 0 180 $X=629920 $Y=733900
X1540 3698 3314 3592 2 1 3658 QDFFRBN $T=643560 850200 1 180 $X=631780 $Y=849820
X1541 3711 622 577 2 1 599 QDFFRBN $T=644800 890520 0 180 $X=633020 $Y=885100
X1542 3674 550 3519 2 1 628 QDFFRBN $T=634260 739320 0 0 $X=634260 $Y=738940
X1543 3718 550 3641 2 1 3670 QDFFRBN $T=646040 749400 0 180 $X=634260 $Y=743980
X1544 3672 3314 3687 2 1 631 QDFFRBN $T=634260 870360 1 0 $X=634260 $Y=864940
X1545 3676 550 3712 2 1 3727 QDFFRBN $T=635500 769560 1 0 $X=635500 $Y=764140
X1546 3677 3314 3657 2 1 616 QDFFRBN $T=635500 830040 0 0 $X=635500 $Y=829660
X1547 610 550 3544 2 1 632 QDFFRBN $T=636120 729240 0 0 $X=636120 $Y=728860
X1548 3730 622 3667 2 1 3661 QDFFRBN $T=651620 880440 1 180 $X=639840 $Y=880060
X1549 3741 622 3644 2 1 3695 QDFFRBN $T=652240 779640 1 180 $X=640460 $Y=779260
X1550 3702 3314 3687 2 1 3689 QDFFRBN $T=641700 880440 1 0 $X=641700 $Y=875020
X1551 3715 3314 3742 2 1 3758 QDFFRBN $T=642940 840120 0 0 $X=642940 $Y=839740
X1552 3710 3314 3742 2 1 3751 QDFFRBN $T=642940 860280 0 0 $X=642940 $Y=859900
X1553 3763 550 3519 2 1 626 QDFFRBN $T=655340 739320 0 180 $X=643560 $Y=733900
X1554 3716 3314 3750 2 1 3709 QDFFRBN $T=643560 809880 1 0 $X=643560 $Y=804460
X1555 3708 3314 3654 2 1 3651 QDFFRBN $T=643560 809880 0 0 $X=643560 $Y=809500
X1556 3717 3314 3742 2 1 3766 QDFFRBN $T=643560 850200 0 0 $X=643560 $Y=849820
X1557 3721 622 3654 2 1 614 QDFFRBN $T=655960 819960 1 180 $X=644180 $Y=819580
X1558 3722 3314 3687 2 1 3588 QDFFRBN $T=645420 870360 0 0 $X=645420 $Y=869980
X1559 3781 550 3641 2 1 3723 QDFFRBN $T=657820 749400 0 180 $X=646040 $Y=743980
X1560 3756 622 3654 2 1 3701 QDFFRBN $T=657820 830040 0 180 $X=646040 $Y=824620
X1561 3733 622 3712 2 1 3754 QDFFRBN $T=647280 769560 1 0 $X=647280 $Y=764140
X1562 3731 622 3644 2 1 2662 QDFFRBN $T=660920 789720 1 180 $X=649140 $Y=789340
X1563 3760 622 3800 2 1 3776 QDFFRBN $T=652860 789720 1 0 $X=652860 $Y=784300
X1564 3768 550 3779 2 1 660 QDFFRBN $T=654720 729240 0 0 $X=654720 $Y=728860
X1565 3774 622 3712 2 1 3780 QDFFRBN $T=655340 779640 1 0 $X=655340 $Y=774220
X1566 3820 550 3712 2 1 647 QDFFRBN $T=668360 759480 0 180 $X=656580 $Y=754060
X1567 3798 622 3797 2 1 3675 QDFFRBN $T=668980 819960 1 180 $X=657200 $Y=819580
X1568 3783 622 3742 2 1 665 QDFFRBN $T=657200 860280 0 0 $X=657200 $Y=859900
X1569 3784 550 3779 2 1 667 QDFFRBN $T=657820 739320 1 0 $X=657820 $Y=733900
X1570 3786 622 3750 2 1 3682 QDFFRBN $T=657820 819960 1 0 $X=657820 $Y=814540
X1571 3788 622 3742 2 1 3560 QDFFRBN $T=658440 850200 0 0 $X=658440 $Y=849820
X1572 3789 622 3742 2 1 3812 QDFFRBN $T=659060 840120 0 0 $X=659060 $Y=839740
X1573 3799 550 3641 2 1 3819 QDFFRBN $T=660300 749400 0 0 $X=660300 $Y=749020
X1574 3804 622 3837 2 1 3849 QDFFRBN $T=660920 880440 0 0 $X=660920 $Y=880060
X1575 3805 622 666 2 1 3726 QDFFRBN $T=660920 900600 1 0 $X=660920 $Y=895180
X1576 3811 622 3750 2 1 3861 QDFFRBN $T=662160 809880 0 0 $X=662160 $Y=809500
X1577 3817 622 3800 2 1 3845 QDFFRBN $T=664020 779640 0 0 $X=664020 $Y=779260
X1578 3824 622 3797 2 1 3865 QDFFRBN $T=665260 830040 1 0 $X=665260 $Y=824620
X1579 3823 550 3864 2 1 3790 QDFFRBN $T=665880 739320 0 0 $X=665880 $Y=738940
X1580 3855 622 3800 2 1 3826 QDFFRBN $T=677660 789720 0 180 $X=665880 $Y=784300
X1581 3840 622 3797 2 1 3284 QDFFRBN $T=669600 830040 0 0 $X=669600 $Y=829660
X1582 3848 622 3837 2 1 693 QDFFRBN $T=671460 880440 1 0 $X=671460 $Y=875020
X1583 3851 550 3864 2 1 694 QDFFRBN $T=672080 739320 1 0 $X=672080 $Y=733900
X1584 3853 622 3837 2 1 3703 QDFFRBN $T=672080 860280 0 0 $X=672080 $Y=859900
X1585 3914 622 3800 2 1 3860 QDFFRBN $T=685100 779640 0 180 $X=673320 $Y=774220
X1586 3863 622 3837 2 1 3814 QDFFRBN $T=673320 870360 0 0 $X=673320 $Y=869980
X1587 3866 622 3837 2 1 3810 QDFFRBN $T=673940 890520 1 0 $X=673940 $Y=885100
X1588 3886 622 3881 2 1 3854 QDFFRBN $T=686960 769560 0 180 $X=675180 $Y=764140
X1589 3899 622 3750 2 1 3831 QDFFRBN $T=687580 809880 0 180 $X=675800 $Y=804460
X1590 3938 622 3797 2 1 3876 QDFFRBN $T=688820 830040 0 180 $X=677040 $Y=824620
X1591 3945 550 3864 2 1 3885 QDFFRBN $T=690680 739320 1 180 $X=678900 $Y=738940
X1592 3908 622 3881 2 1 710 QDFFRBN $T=682000 789720 1 0 $X=682000 $Y=784300
X1593 3909 622 3887 2 1 3961 QDFFRBN $T=682000 799800 0 0 $X=682000 $Y=799420
X1594 3882 622 3955 2 1 3728 QDFFRBN $T=682620 840120 0 0 $X=682620 $Y=839740
X1595 3915 622 3887 2 1 3953 QDFFRBN $T=683240 809880 0 0 $X=683240 $Y=809500
X1596 3927 550 3864 2 1 3963 QDFFRBN $T=685720 739320 1 0 $X=685720 $Y=733900
X1597 3984 622 3951 2 1 3932 QDFFRBN $T=698120 860280 1 180 $X=686340 $Y=859900
X1598 3990 622 3881 2 1 3929 QDFFRBN $T=700600 769560 0 180 $X=688820 $Y=764140
X1599 4005 622 3797 2 1 3944 QDFFRBN $T=700600 830040 0 180 $X=688820 $Y=824620
X1600 4010 550 3864 2 1 3952 QDFFRBN $T=703080 739320 1 180 $X=691300 $Y=738940
X1601 3968 622 725 2 1 4008 QDFFRBN $T=692540 900600 1 0 $X=692540 $Y=895180
X1602 4032 622 3881 2 1 3977 QDFFRBN $T=706180 779640 1 180 $X=694400 $Y=779260
X1603 3993 622 3955 2 1 703 QDFFRBN $T=706800 840120 1 180 $X=695020 $Y=839740
X1604 4064 622 4007 2 1 3987 QDFFRBN $T=708040 799800 1 180 $X=696260 $Y=799420
X1605 4028 622 4007 2 1 3917 QDFFRBN $T=709900 789720 1 180 $X=698120 $Y=789340
X1606 4059 550 719 2 1 4015 QDFFRBN $T=712380 739320 0 180 $X=700600 $Y=733900
X1607 4021 622 3951 2 1 4056 QDFFRBN $T=700600 860280 0 0 $X=700600 $Y=859900
X1608 4073 550 3779 2 1 4023 QDFFRBN $T=713000 749400 0 180 $X=701220 $Y=743980
X1609 4090 622 725 2 1 3985 QDFFRBN $T=713620 890520 0 180 $X=701840 $Y=885100
X1610 4045 622 4007 2 1 4058 QDFFRBN $T=704320 789720 1 0 $X=704320 $Y=784300
X1611 4096 622 4139 2 1 4091 QDFFRBN $T=713000 819960 0 0 $X=713000 $Y=819580
X1612 4153 760 4123 2 1 4103 QDFFRBN $T=725400 860280 1 180 $X=713620 $Y=859900
X1613 4154 622 751 2 1 4070 QDFFRBN $T=725400 890520 0 180 $X=713620 $Y=885100
X1614 4108 4151 4007 2 1 4037 QDFFRBN $T=726020 799800 0 180 $X=714240 $Y=794380
X1615 4087 761 4129 2 1 744 QDFFRBN $T=726640 749400 0 180 $X=714860 $Y=743980
X1616 4116 622 4139 2 1 4077 QDFFRBN $T=714860 809880 1 0 $X=714860 $Y=804460
X1617 4134 761 755 2 1 4113 QDFFRBN $T=727260 739320 0 180 $X=715480 $Y=733900
X1618 4143 4151 4129 2 1 4095 QDFFRBN $T=727260 759480 1 180 $X=715480 $Y=759100
X1619 4128 4151 4129 2 1 4122 QDFFRBN $T=729120 759480 0 180 $X=717340 $Y=754060
X1620 4106 4151 4129 2 1 736 QDFFRBN $T=729120 779640 1 180 $X=717340 $Y=779260
X1621 4114 4151 4139 2 1 4082 QDFFRBN $T=729120 799800 1 180 $X=717340 $Y=799420
X1622 4166 760 4123 2 1 4068 QDFFRBN $T=729120 870360 0 180 $X=717340 $Y=864940
X1623 4168 4151 4139 2 1 4111 QDFFRBN $T=729740 819960 0 180 $X=717960 $Y=814540
X1624 4105 760 751 2 1 4072 QDFFRBN $T=729740 900600 0 180 $X=717960 $Y=895180
X1625 4163 4151 4129 2 1 742 QDFFRBN $T=730980 769560 0 180 $X=719200 $Y=764140
X1626 4147 761 755 2 1 774 QDFFRBN $T=721680 739320 0 0 $X=721680 $Y=738940
X1627 4156 4151 4192 2 1 4117 QDFFRBN $T=724780 830040 0 0 $X=724780 $Y=829660
X1628 4216 760 751 2 1 770 QDFFRBN $T=739040 890520 0 180 $X=727260 $Y=885100
X1629 4169 760 4123 2 1 4249 QDFFRBN $T=727880 880440 0 0 $X=727880 $Y=880060
X1630 4171 4151 4193 2 1 794 QDFFRBN $T=728500 809880 1 0 $X=728500 $Y=804460
X1631 4172 760 4123 2 1 4214 QDFFRBN $T=728500 880440 1 0 $X=728500 $Y=875020
X1632 810 4151 4224 2 1 4191 QDFFRBN $T=746480 769560 0 180 $X=734700 $Y=764140
X1633 4207 761 808 2 1 816 QDFFRBN $T=735320 729240 0 0 $X=735320 $Y=728860
X1634 4239 4151 4192 2 1 4206 QDFFRBN $T=748340 830040 1 180 $X=736560 $Y=829660
X1635 4286 4151 4193 2 1 4223 QDFFRBN $T=752060 809880 0 180 $X=740280 $Y=804460
X1636 4245 760 4192 2 1 4184 QDFFRBN $T=752060 840120 0 180 $X=740280 $Y=834700
X1637 4283 760 4192 2 1 4228 QDFFRBN $T=755780 850200 1 180 $X=744000 $Y=849820
X1638 4269 4151 4304 2 1 4227 QDFFRBN $T=745240 830040 1 0 $X=745240 $Y=824620
X1639 4261 760 751 2 1 4187 QDFFRBN $T=758260 890520 0 180 $X=746480 $Y=885100
X1640 4262 760 822 2 1 796 QDFFRBN $T=758260 900600 0 180 $X=746480 $Y=895180
X1641 4274 761 808 2 1 4307 QDFFRBN $T=747100 729240 1 0 $X=747100 $Y=723820
X1642 4254 4151 4304 2 1 4217 QDFFRBN $T=747720 819960 0 0 $X=747720 $Y=819580
X1643 4277 760 4317 2 1 4247 QDFFRBN $T=747720 880440 1 0 $X=747720 $Y=875020
X1644 4291 760 4330 2 1 4231 QDFFRBN $T=750200 870360 0 0 $X=750200 $Y=869980
X1645 4342 4151 4192 2 1 4200 QDFFRBN $T=762600 830040 1 180 $X=750820 $Y=829660
X1646 4297 4151 4193 2 1 844 QDFFRBN $T=752060 809880 1 0 $X=752060 $Y=804460
X1647 4298 4151 4304 2 1 845 QDFFRBN $T=752060 819960 1 0 $X=752060 $Y=814540
X1648 4301 760 4330 2 1 4369 QDFFRBN $T=752680 860280 1 0 $X=752680 $Y=854860
X1649 4305 760 4304 2 1 4325 QDFFRBN $T=753300 850200 1 0 $X=753300 $Y=844780
X1650 4296 760 4123 2 1 807 QDFFRBN $T=765700 860280 1 180 $X=753920 $Y=859900
X1651 4319 4151 4193 2 1 4368 QDFFRBN $T=755780 789720 0 0 $X=755780 $Y=789340
X1652 4320 4151 4193 2 1 853 QDFFRBN $T=755780 799800 1 0 $X=755780 $Y=794380
X1653 4321 4151 4193 2 1 852 QDFFRBN $T=755780 799800 0 0 $X=755780 $Y=799420
X1654 4333 4151 4304 2 1 4390 QDFFRBN $T=758880 830040 1 0 $X=758880 $Y=824620
X1655 4339 4151 4382 2 1 4401 QDFFRBN $T=760120 819960 0 0 $X=760120 $Y=819580
X1656 4340 760 822 2 1 4392 QDFFRBN $T=760120 900600 1 0 $X=760120 $Y=895180
X1657 4354 760 4317 2 1 4358 QDFFRBN $T=762600 880440 1 0 $X=762600 $Y=875020
X1658 4364 760 4330 2 1 4341 QDFFRBN $T=765700 870360 1 0 $X=765700 $Y=864940
X1659 4375 760 4317 2 1 4258 QDFFRBN $T=766940 870360 0 0 $X=766940 $Y=869980
X1660 4469 761 4433 2 1 864 QDFFRBN $T=784920 759480 1 180 $X=773140 $Y=759100
X1661 4476 761 4433 2 1 4416 QDFFRBN $T=785540 749400 1 180 $X=773760 $Y=749020
X1662 4417 4151 4462 2 1 4443 QDFFRBN $T=773760 809880 0 0 $X=773760 $Y=809500
X1663 4465 760 4382 2 1 4438 QDFFRBN $T=788020 840120 1 180 $X=776240 $Y=839740
X1664 4445 760 4475 2 1 854 QDFFRBN $T=776860 890520 1 0 $X=776860 $Y=885100
X1665 4442 4151 4467 2 1 889 QDFFRBN $T=779340 769560 0 0 $X=779340 $Y=769180
X1666 4459 760 4317 2 1 898 QDFFRBN $T=780580 870360 0 0 $X=780580 $Y=869980
X1667 4533 4151 4462 2 1 4468 QDFFRBN $T=794840 830040 1 180 $X=783060 $Y=829660
X1668 4471 760 4475 2 1 4452 QDFFRBN $T=783060 900600 1 0 $X=783060 $Y=895180
X1669 4542 760 4330 2 1 4478 QDFFRBN $T=796080 850200 0 180 $X=784300 $Y=844780
X1670 4552 761 4433 2 1 4486 QDFFRBN $T=797320 739320 1 180 $X=785540 $Y=738940
X1671 4557 761 4433 2 1 884 QDFFRBN $T=797940 729240 1 180 $X=786160 $Y=728860
X1672 4494 4151 4462 2 1 4513 QDFFRBN $T=786160 809880 0 0 $X=786160 $Y=809500
X1673 4573 761 4433 2 1 894 QDFFRBN $T=799800 729240 0 180 $X=788020 $Y=723820
X1674 4493 4151 4462 2 1 4362 QDFFRBN $T=788020 830040 1 0 $X=788020 $Y=824620
X1675 4515 4151 4467 2 1 4504 QDFFRBN $T=800420 779640 1 180 $X=788640 $Y=779260
X1676 4549 760 4461 2 1 896 QDFFRBN $T=800420 880440 0 180 $X=788640 $Y=875020
X1677 4562 4151 4433 2 1 4511 QDFFRBN $T=801040 759480 0 180 $X=789260 $Y=754060
X1678 4558 4151 4467 2 1 902 QDFFRBN $T=806000 769560 1 180 $X=794220 $Y=769180
X1679 4526 4151 4576 2 1 4335 QDFFRBN $T=794840 809880 1 0 $X=794840 $Y=804460
X1680 4559 4151 4576 2 1 4616 QDFFRBN $T=796080 789720 1 0 $X=796080 $Y=784300
X1681 4569 760 4461 2 1 4536 QDFFRBN $T=809100 880440 1 180 $X=797320 $Y=880060
X1682 4633 4151 4582 2 1 4510 QDFFRBN $T=809720 809880 1 180 $X=797940 $Y=809500
X1683 4634 760 4583 2 1 4568 QDFFRBN $T=809720 850200 0 180 $X=797940 $Y=844780
X1684 4609 4151 4462 2 1 4501 QDFFRBN $T=812200 830040 0 180 $X=800420 $Y=824620
X1685 4586 4151 4639 2 1 4597 QDFFRBN $T=801040 759480 1 0 $X=801040 $Y=754060
X1686 4652 4151 4462 2 1 914 QDFFRBN $T=812820 819960 0 180 $X=801040 $Y=814540
X1687 4592 761 4639 2 1 4588 QDFFRBN $T=801660 749400 1 0 $X=801660 $Y=743980
X1688 4653 760 4556 2 1 4601 QDFFRBN $T=814680 880440 0 180 $X=802900 $Y=875020
X1689 4561 760 4556 2 1 918 QDFFRBN $T=804140 900600 1 0 $X=804140 $Y=895180
X1690 4673 4151 4576 2 1 4617 QDFFRBN $T=818400 809880 0 180 $X=806620 $Y=804460
X1691 4661 933 4639 2 1 920 QDFFRBN $T=819020 739320 1 180 $X=807240 $Y=738940
X1692 4614 4151 4639 2 1 4571 QDFFRBN $T=809100 769560 0 0 $X=809100 $Y=769180
X1693 4640 4151 4583 2 1 4670 QDFFRBN $T=809100 830040 0 0 $X=809100 $Y=829660
X1694 4698 937 912 2 1 919 QDFFRBN $T=820880 890520 1 180 $X=809100 $Y=890140
X1695 4690 4151 4582 2 1 4643 QDFFRBN $T=823360 789720 0 180 $X=811580 $Y=784300
X1696 4715 760 4583 2 1 4567 QDFFRBN $T=823360 840120 1 180 $X=811580 $Y=839740
X1697 4678 933 4639 2 1 4744 QDFFRBN $T=815920 759480 0 0 $X=815920 $Y=759100
X1698 4682 933 4728 2 1 4723 QDFFRBN $T=816540 749400 0 0 $X=816540 $Y=749020
X1699 4745 4151 4582 2 1 4629 QDFFRBN $T=830180 789720 1 180 $X=818400 $Y=789340
X1700 4765 4151 4582 2 1 4691 QDFFRBN $T=830180 809880 0 180 $X=818400 $Y=804460
X1701 4693 4151 4741 2 1 4565 QDFFRBN $T=818400 809880 0 0 $X=818400 $Y=809500
X1702 4696 4151 4688 2 1 4761 QDFFRBN $T=819020 830040 1 0 $X=819020 $Y=824620
X1703 4697 937 4556 2 1 4763 QDFFRBN $T=819020 890520 1 0 $X=819020 $Y=885100
X1704 4709 933 4728 2 1 4768 QDFFRBN $T=820880 739320 1 0 $X=820880 $Y=733900
X1705 4767 933 4728 2 1 4711 QDFFRBN $T=833280 739320 1 180 $X=821500 $Y=738940
X1706 4718 4151 4741 2 1 4554 QDFFRBN $T=822120 819960 1 0 $X=822120 $Y=814540
X1707 4729 4151 4688 2 1 4522 QDFFRBN $T=823980 819960 0 0 $X=823980 $Y=819580
X1708 4733 4151 4725 2 1 4779 QDFFRBN $T=825220 769560 0 0 $X=825220 $Y=769180
X1709 4742 760 4688 2 1 4735 QDFFRBN $T=826460 850200 1 0 $X=826460 $Y=844780
X1710 4797 937 4712 2 1 4737 QDFFRBN $T=838860 860280 1 180 $X=827080 $Y=859900
X1711 4807 937 912 2 1 4749 QDFFRBN $T=839480 900600 0 180 $X=827700 $Y=895180
X1712 4727 937 4712 2 1 4730 QDFFRBN $T=845060 860280 0 180 $X=833280 $Y=854860
X1713 4799 933 4806 2 1 4817 QDFFRBN $T=836380 749400 1 0 $X=836380 $Y=743980
X1714 4861 933 4806 2 1 4808 QDFFRBN $T=850020 749400 1 180 $X=838240 $Y=749020
X1715 4809 4151 4847 2 1 4848 QDFFRBN $T=838240 769560 1 0 $X=838240 $Y=764140
X1716 4838 937 4556 2 1 4598 QDFFRBN $T=850020 890520 0 180 $X=838240 $Y=885100
X1717 4811 4151 4741 2 1 4842 QDFFRBN $T=838860 809880 1 0 $X=838860 $Y=804460
X1718 4844 4850 4725 2 1 4795 QDFFRBN $T=851260 779640 0 180 $X=839480 $Y=774220
X1719 4862 933 968 2 1 4818 QDFFRBN $T=852500 729240 1 180 $X=840720 $Y=728860
X1720 4793 937 4852 2 1 4774 QDFFRBN $T=840720 830040 1 0 $X=840720 $Y=824620
X1721 4823 937 4852 2 1 4812 QDFFRBN $T=840720 840120 0 0 $X=840720 $Y=839740
X1722 4832 937 972 2 1 4798 QDFFRBN $T=842580 900600 1 0 $X=842580 $Y=895180
X1723 4869 937 4839 2 1 4313 QDFFRBN $T=854980 870360 1 180 $X=843200 $Y=869980
X1724 4868 4850 4852 2 1 4611 QDFFRBN $T=856220 830040 1 180 $X=844440 $Y=829660
X1725 4855 4850 4900 2 1 4637 QDFFRBN $T=846920 799800 1 0 $X=846920 $Y=794380
X1726 4860 937 4911 2 1 4930 QDFFRBN $T=848780 890520 0 0 $X=848780 $Y=890140
X1727 4865 4850 4847 2 1 4926 QDFFRBN $T=849400 779640 0 0 $X=849400 $Y=779260
X1728 4880 4850 4741 2 1 4875 QDFFRBN $T=851880 809880 0 0 $X=851880 $Y=809500
X1729 4886 4850 4900 2 1 4943 QDFFRBN $T=852500 789720 0 0 $X=852500 $Y=789340
X1730 4894 4850 4847 2 1 984 QDFFRBN $T=853120 779640 1 0 $X=853120 $Y=774220
X1731 4896 4850 4741 2 1 4906 QDFFRBN $T=853740 809880 1 0 $X=853740 $Y=804460
X1732 977 933 968 2 1 4959 QDFFRBN $T=854360 729240 0 0 $X=854360 $Y=728860
X1733 4864 4850 4919 2 1 4858 QDFFRBN $T=868000 819960 1 180 $X=856220 $Y=819580
X1734 4944 4850 4839 2 1 4907 QDFFRBN $T=868000 850200 0 180 $X=856220 $Y=844780
X1735 4954 4850 4919 2 1 4757 QDFFRBN $T=868620 830040 0 180 $X=856840 $Y=824620
X1736 4905 4850 4948 2 1 4934 QDFFRBN $T=857460 759480 0 0 $X=857460 $Y=759100
X1737 4937 937 4927 2 1 969 QDFFRBN $T=869240 870360 1 180 $X=857460 $Y=869980
X1738 4962 4850 4919 2 1 4671 QDFFRBN $T=869860 830040 1 180 $X=858080 $Y=829660
X1739 4917 937 980 2 1 4831 QDFFRBN $T=858080 900600 1 0 $X=858080 $Y=895180
X1740 4921 937 4839 2 1 4942 QDFFRBN $T=859320 860280 0 0 $X=859320 $Y=859900
X1741 4913 937 4911 2 1 4825 QDFFRBN $T=871100 880440 1 180 $X=859320 $Y=880060
X1742 4940 933 968 2 1 4898 QDFFRBN $T=871720 739320 0 180 $X=859940 $Y=733900
X1743 4989 4850 4919 2 1 4936 QDFFRBN $T=874200 840120 1 180 $X=862420 $Y=839740
X1744 5005 4850 4847 2 1 4938 QDFFRBN $T=874820 779640 1 180 $X=863040 $Y=779260
X1745 4951 937 4927 2 1 5000 QDFFRBN $T=865520 880440 1 0 $X=865520 $Y=875020
X1746 4966 4850 4900 2 1 4956 QDFFRBN $T=868620 819960 1 0 $X=868620 $Y=814540
X1747 4967 4850 4948 2 1 4994 QDFFRBN $T=869240 759480 1 0 $X=869240 $Y=754060
X1748 4971 4850 4948 2 1 5004 QDFFRBN $T=870480 769560 1 0 $X=870480 $Y=764140
X1749 4960 4850 5020 2 1 4958 QDFFRBN $T=870480 799800 0 0 $X=870480 $Y=799420
X1750 4985 937 4927 2 1 5046 QDFFRBN $T=871720 860280 0 0 $X=871720 $Y=859900
X1751 4986 937 990 2 1 4973 QDFFRBN $T=871720 880440 0 0 $X=871720 $Y=880060
X1752 4988 4850 5021 2 1 5022 QDFFRBN $T=872340 830040 0 0 $X=872340 $Y=829660
X1753 4987 933 5034 2 1 5015 QDFFRBN $T=872960 729240 0 0 $X=872960 $Y=728860
X1754 5051 937 4927 2 1 4993 QDFFRBN $T=884740 870360 0 180 $X=872960 $Y=864940
X1755 5011 4850 5020 2 1 4980 QDFFRBN $T=887220 809880 1 180 $X=875440 $Y=809500
X1756 5063 4850 5042 2 1 5023 QDFFRBN $T=890940 769560 1 180 $X=879160 $Y=769180
X1757 1008 933 5034 2 1 1021 QDFFRBN $T=881640 729240 1 0 $X=881640 $Y=723820
X1758 5107 4850 4948 2 1 1007 QDFFRBN $T=894660 759480 0 180 $X=882880 $Y=754060
X1759 5050 4850 5020 2 1 5120 QDFFRBN $T=882880 809880 1 0 $X=882880 $Y=804460
X1760 5109 937 4911 2 1 5047 QDFFRBN $T=894660 880440 0 180 $X=882880 $Y=875020
X1761 5054 4850 5020 2 1 5006 QDFFRBN $T=883500 799800 0 0 $X=883500 $Y=799420
X1762 5097 933 5034 2 1 5069 QDFFRBN $T=898380 739320 1 180 $X=886600 $Y=738940
X1763 5123 933 5034 2 1 1013 QDFFRBN $T=899000 729240 1 180 $X=887220 $Y=728860
X1764 5082 4850 5042 2 1 5153 QDFFRBN $T=887840 779640 1 0 $X=887840 $Y=774220
X1765 5126 937 5021 2 1 5083 QDFFRBN $T=900240 850200 1 180 $X=888460 $Y=849820
X1766 5135 937 5101 2 1 5084 QDFFRBN $T=900240 870360 0 180 $X=888460 $Y=864940
X1767 5133 937 990 2 1 5048 QDFFRBN $T=902100 890520 0 180 $X=890320 $Y=885100
X1768 5085 937 990 2 1 997 QDFFRBN $T=902100 900600 0 180 $X=890320 $Y=895180
X1769 5104 4850 5117 2 1 5165 QDFFRBN $T=891560 819960 0 0 $X=891560 $Y=819580
X1770 5094 937 5021 2 1 5065 QDFFRBN $T=904580 840120 1 180 $X=892800 $Y=839740
X1771 5110 937 990 2 1 5147 QDFFRBN $T=892800 880440 0 0 $X=892800 $Y=880060
X1772 5161 4850 4948 2 1 1016 QDFFRBN $T=905200 769560 1 180 $X=893420 $Y=769180
X1773 5143 4850 5042 2 1 5115 QDFFRBN $T=905820 779640 1 180 $X=894040 $Y=779260
X1774 5158 4850 5034 2 1 5087 QDFFRBN $T=908920 759480 0 180 $X=897140 $Y=754060
X1775 5099 4850 5181 2 1 1010 QDFFRBN $T=897140 799800 0 0 $X=897140 $Y=799420
X1776 5184 4850 5117 2 1 5155 QDFFRBN $T=913260 830040 0 180 $X=901480 $Y=824620
X1777 5213 4850 5117 2 1 5132 QDFFRBN $T=913260 830040 1 180 $X=901480 $Y=829660
X1778 5218 937 5101 2 1 5170 QDFFRBN $T=915740 880440 0 180 $X=903960 $Y=875020
X1779 5206 937 5191 2 1 5142 QDFFRBN $T=915740 890520 0 180 $X=903960 $Y=885100
X1780 5222 4850 5042 2 1 5116 QDFFRBN $T=918220 779640 1 180 $X=906440 $Y=779260
X1781 5171 1043 1036 2 1 5149 QDFFRBN $T=918840 729240 0 180 $X=907060 $Y=723820
X1782 5198 4850 5181 2 1 5134 QDFFRBN $T=919460 789720 1 180 $X=907680 $Y=789340
X1783 5197 4850 5225 2 1 5241 QDFFRBN $T=908300 759480 0 0 $X=908300 $Y=759100
X1784 5167 4850 5226 2 1 5144 QDFFRBN $T=908300 840120 1 0 $X=908300 $Y=834700
X1785 5174 937 5227 2 1 4969 QDFFRBN $T=908300 860280 1 0 $X=908300 $Y=854860
X1786 5200 4850 5225 2 1 5235 QDFFRBN $T=908920 779640 1 0 $X=908920 $Y=774220
X1787 5229 4850 5181 2 1 5202 QDFFRBN $T=921320 799800 0 180 $X=909540 $Y=794380
X1788 5196 1045 5191 2 1 1032 QDFFRBN $T=921320 890520 1 180 $X=909540 $Y=890140
X1789 5192 1043 1036 2 1 5160 QDFFRBN $T=921940 729240 1 180 $X=910160 $Y=728860
X1790 5201 1043 1036 2 1 5140 QDFFRBN $T=923180 739320 1 180 $X=911400 $Y=738940
X1791 5199 937 5227 2 1 5166 QDFFRBN $T=912020 850200 1 0 $X=912020 $Y=844780
X1792 5214 4850 1036 2 1 5265 QDFFRBN $T=913260 749400 1 0 $X=913260 $Y=743980
X1793 5219 937 5101 2 1 5264 QDFFRBN $T=913880 880440 0 0 $X=913880 $Y=880060
X1794 5228 4850 5225 2 1 5268 QDFFRBN $T=915740 759480 1 0 $X=915740 $Y=754060
X1795 5223 937 5101 2 1 5270 QDFFRBN $T=915740 870360 0 0 $X=915740 $Y=869980
X1796 5224 937 5101 2 1 1047 QDFFRBN $T=915740 880440 1 0 $X=915740 $Y=875020
X1797 5230 4850 5242 2 1 5299 QDFFRBN $T=916360 830040 1 0 $X=916360 $Y=824620
X1798 5236 4850 5253 2 1 5283 QDFFRBN $T=918840 799800 0 0 $X=918840 $Y=799420
X1799 5238 4850 5253 2 1 5275 QDFFRBN $T=919460 789720 1 0 $X=919460 $Y=784300
X1800 5306 4850 5253 2 1 5237 QDFFRBN $T=931240 789720 1 180 $X=919460 $Y=789340
X1801 5240 1045 1044 2 1 1050 QDFFRBN $T=919460 900600 1 0 $X=919460 $Y=895180
X1802 5246 4850 5225 2 1 5310 QDFFRBN $T=920700 759480 0 0 $X=920700 $Y=759100
X1803 5249 1043 1049 2 1 5255 QDFFRBN $T=921320 729240 1 0 $X=921320 $Y=723820
X1804 5251 1045 5191 2 1 5305 QDFFRBN $T=921320 890520 0 0 $X=921320 $Y=890140
X1805 5254 937 5194 2 1 5216 QDFFRBN $T=922560 850200 0 0 $X=922560 $Y=849820
X1806 5258 4850 5242 2 1 5301 QDFFRBN $T=923180 819960 1 0 $X=923180 $Y=814540
X1807 5239 5317 5253 2 1 5193 QDFFRBN $T=935580 809880 1 180 $X=923800 $Y=809500
X1808 5271 1043 5294 2 1 5342 QDFFRBN $T=926900 749400 1 0 $X=926900 $Y=743980
X1809 5300 1043 1049 2 1 5371 QDFFRBN $T=930620 739320 1 0 $X=930620 $Y=733900
X1810 5314 4850 5361 2 1 5377 QDFFRBN $T=931860 769560 0 0 $X=931860 $Y=769180
X1811 5315 5317 5337 2 1 5372 QDFFRBN $T=931860 799800 0 0 $X=931860 $Y=799420
X1812 5327 4850 5361 2 1 5358 QDFFRBN $T=933720 789720 1 0 $X=933720 $Y=784300
X1813 5389 5317 5242 2 1 5329 QDFFRBN $T=946120 819960 1 180 $X=934340 $Y=819580
X1814 5334 937 5194 2 1 5360 QDFFRBN $T=934960 850200 0 0 $X=934960 $Y=849820
X1815 5336 1045 5384 2 1 5400 QDFFRBN $T=935580 870360 0 0 $X=935580 $Y=869980
X1816 5340 1045 5384 2 1 1068 QDFFRBN $T=936820 890520 1 0 $X=936820 $Y=885100
X1817 5343 5317 5337 2 1 5321 QDFFRBN $T=937440 809880 0 0 $X=937440 $Y=809500
X1818 5429 5317 5226 2 1 5347 QDFFRBN $T=949840 830040 0 180 $X=938060 $Y=824620
X1819 5368 1043 5294 2 1 5405 QDFFRBN $T=940540 749400 1 0 $X=940540 $Y=743980
X1820 5402 1045 1070 2 1 1066 QDFFRBN $T=954180 900600 0 180 $X=942400 $Y=895180
X1821 5423 1045 5384 2 1 5401 QDFFRBN $T=958520 880440 1 180 $X=946740 $Y=880060
X1822 5414 4850 5361 2 1 5481 QDFFRBN $T=947360 789720 1 0 $X=947360 $Y=784300
X1823 5430 5317 5194 2 1 5479 QDFFRBN $T=949840 860280 0 0 $X=949840 $Y=859900
X1824 5489 5317 5337 2 1 5432 QDFFRBN $T=962240 809880 1 180 $X=950460 $Y=809500
X1825 5466 5317 5361 2 1 1072 QDFFRBN $T=964100 799800 0 180 $X=952320 $Y=794380
X1826 5464 5317 5460 2 1 5410 QDFFRBN $T=964100 840120 0 180 $X=952320 $Y=834700
X1827 5433 5317 5194 2 1 5472 QDFFRBN $T=952320 860280 1 0 $X=952320 $Y=854860
X1828 5443 1045 1070 2 1 1079 QDFFRBN $T=952940 890520 0 0 $X=952940 $Y=890140
X1829 5477 5317 5294 2 1 5442 QDFFRBN $T=965960 749400 0 180 $X=954180 $Y=743980
X1830 5467 5317 5384 2 1 5457 QDFFRBN $T=956040 850200 0 0 $X=956040 $Y=849820
X1831 5507 5317 5452 2 1 5469 QDFFRBN $T=968440 779640 0 180 $X=956660 $Y=774220
X1832 5506 1043 1049 2 1 5474 QDFFRBN $T=969060 729240 1 180 $X=957280 $Y=728860
X1833 5517 5317 5361 2 1 5444 QDFFRBN $T=970300 789720 1 180 $X=958520 $Y=789340
X1834 5485 5317 5452 2 1 5550 QDFFRBN $T=959760 769560 1 0 $X=959760 $Y=764140
X1835 5520 5317 5294 2 1 5456 QDFFRBN $T=972160 749400 1 180 $X=960380 $Y=749020
X1836 5516 5317 5564 2 1 5551 QDFFRBN $T=965340 799800 0 0 $X=965340 $Y=799420
X1837 5505 5317 5460 2 1 5465 QDFFRBN $T=965960 840120 1 0 $X=965960 $Y=834700
X1838 5570 5317 5454 2 1 5524 QDFFRBN $T=978980 819960 0 180 $X=967200 $Y=814540
X1839 5584 5317 5460 2 1 5525 QDFFRBN $T=978980 830040 0 180 $X=967200 $Y=824620
X1840 5531 1045 5536 2 1 5543 QDFFRBN $T=967200 890520 0 0 $X=967200 $Y=890140
X1841 5533 5317 5384 2 1 5573 QDFFRBN $T=968440 860280 1 0 $X=968440 $Y=854860
X1842 5611 5317 5454 2 1 5513 QDFFRBN $T=981460 809880 0 180 $X=969680 $Y=804460
X1843 5561 1043 1049 2 1 5534 QDFFRBN $T=982080 729240 1 180 $X=970300 $Y=728860
X1844 5571 5317 5384 2 1 5547 QDFFRBN $T=983940 850200 1 180 $X=972160 $Y=849820
X1845 5566 5317 5608 2 1 5530 QDFFRBN $T=972780 789720 1 0 $X=972780 $Y=784300
X1846 5592 1045 5536 2 1 5540 QDFFRBN $T=985180 880440 1 180 $X=973400 $Y=880060
X1847 5593 5317 5608 2 1 5542 QDFFRBN $T=990140 789720 1 180 $X=978360 $Y=789340
X1848 5585 5317 5640 2 1 5637 QDFFRBN $T=978980 860280 0 0 $X=978980 $Y=859900
X1849 5633 1045 5536 2 1 5582 QDFFRBN $T=992620 870360 0 180 $X=980840 $Y=864940
X1850 5622 5317 5640 2 1 5658 QDFFRBN $T=981460 860280 1 0 $X=981460 $Y=854860
X1851 5615 5317 5568 2 1 5580 QDFFRBN $T=994480 769560 0 180 $X=982700 $Y=764140
X1852 5627 5317 5639 2 1 5673 QDFFRBN $T=982700 809880 1 0 $X=982700 $Y=804460
X1853 5629 1045 1108 2 1 5662 QDFFRBN $T=982700 890520 1 0 $X=982700 $Y=885100
X1854 5631 1045 1107 2 1 1112 QDFFRBN $T=983320 900600 1 0 $X=983320 $Y=895180
X1855 5614 1043 1109 2 1 1100 QDFFRBN $T=983940 729240 0 0 $X=983940 $Y=728860
X1856 5624 1043 5568 2 1 5588 QDFFRBN $T=995720 749400 0 180 $X=983940 $Y=743980
X1857 5630 5317 5639 2 1 5599 QDFFRBN $T=995720 830040 0 180 $X=983940 $Y=824620
X1858 5634 5317 5651 2 1 5579 QDFFRBN $T=983940 850200 1 0 $X=983940 $Y=844780
X1859 5625 1043 5568 2 1 5518 QDFFRBN $T=996340 749400 1 180 $X=984560 $Y=749020
X1860 5646 1043 5568 2 1 5598 QDFFRBN $T=996340 759480 0 180 $X=984560 $Y=754060
X1861 5635 5317 5608 2 1 5652 QDFFRBN $T=984560 799800 1 0 $X=984560 $Y=794380
X1862 5632 5317 5639 2 1 5603 QDFFRBN $T=997580 830040 1 180 $X=985800 $Y=829660
X1863 5642 5317 5651 2 1 5607 QDFFRBN $T=986420 840120 0 0 $X=986420 $Y=839740
X1864 5643 5317 5608 2 1 5682 QDFFRBN $T=987040 789720 1 0 $X=987040 $Y=784300
X1865 5676 1045 1108 2 1 5641 QDFFRBN $T=998820 880440 1 180 $X=987040 $Y=880060
X1866 5696 1045 5640 2 1 5645 QDFFRBN $T=1000680 880440 0 180 $X=988900 $Y=875020
X1867 5725 5317 5568 2 1 5650 QDFFRBN $T=1002540 759480 1 180 $X=990760 $Y=759100
X1868 5753 5317 5657 2 1 1111 QDFFRBN $T=1005640 850200 1 180 $X=993860 $Y=849820
X1869 5699 1043 1109 2 1 5656 QDFFRBN $T=1008740 729240 1 180 $X=996960 $Y=728860
X1870 5752 5317 5640 2 1 5679 QDFFRBN $T=1009360 850200 0 180 $X=997580 $Y=844780
X1871 5743 5765 5608 2 1 5693 QDFFRBN $T=1011220 799800 0 180 $X=999440 $Y=794380
X1872 5710 5317 5766 2 1 5737 QDFFRBN $T=1000680 830040 1 0 $X=1000680 $Y=824620
X1873 5721 5317 5766 2 1 5744 QDFFRBN $T=1001920 809880 1 0 $X=1001920 $Y=804460
X1874 5718 5317 5766 2 1 5741 QDFFRBN $T=1001920 819960 0 0 $X=1001920 $Y=819580
X1875 5722 1043 1135 2 1 5789 QDFFRBN $T=1002540 749400 1 0 $X=1002540 $Y=743980
X1876 5738 1045 5774 2 1 1128 QDFFRBN $T=1004400 890520 1 0 $X=1004400 $Y=885100
X1877 1131 1043 1135 2 1 1142 QDFFRBN $T=1006260 729240 1 0 $X=1006260 $Y=723820
X1878 5751 1043 1135 2 1 5777 QDFFRBN $T=1006260 739320 1 0 $X=1006260 $Y=733900
X1879 5810 5317 5651 2 1 5756 QDFFRBN $T=1018660 840120 1 180 $X=1006880 $Y=839740
X1880 5788 1146 5774 2 1 5757 QDFFRBN $T=1018660 870360 0 180 $X=1006880 $Y=864940
X1881 5780 5317 5819 2 1 5812 QDFFRBN $T=1011220 759480 0 0 $X=1011220 $Y=759100
X1882 5783 5317 5774 2 1 5786 QDFFRBN $T=1011840 860280 1 0 $X=1011840 $Y=854860
X1883 5792 5317 5819 2 1 5692 QDFFRBN $T=1013080 779640 1 0 $X=1013080 $Y=774220
X1884 5793 5765 5805 2 1 5848 QDFFRBN $T=1013700 799800 1 0 $X=1013700 $Y=794380
X1885 5795 5765 5805 2 1 5854 QDFFRBN $T=1014320 799800 0 0 $X=1014320 $Y=799420
X1886 5808 1043 1135 2 1 1155 QDFFRBN $T=1016800 729240 0 0 $X=1016800 $Y=728860
X1887 5809 5765 5805 2 1 5847 QDFFRBN $T=1016800 789720 0 0 $X=1016800 $Y=789340
X1888 5811 1045 5774 2 1 5790 QDFFRBN $T=1017420 890520 1 0 $X=1017420 $Y=885100
X1889 5818 5317 5657 2 1 5872 QDFFRBN $T=1018660 830040 0 0 $X=1018660 $Y=829660
X1890 5822 1146 5774 2 1 5884 QDFFRBN $T=1019280 860280 0 0 $X=1019280 $Y=859900
X1891 5862 5765 5657 2 1 5821 QDFFRBN $T=1031680 840120 1 180 $X=1019900 $Y=839740
X1892 5825 1043 5853 2 1 5846 QDFFRBN $T=1020520 739320 1 0 $X=1020520 $Y=733900
X1893 5824 1146 5774 2 1 5879 QDFFRBN $T=1020520 870360 1 0 $X=1020520 $Y=864940
X1894 5837 5317 5819 2 1 5909 QDFFRBN $T=1023000 759480 0 0 $X=1023000 $Y=759100
X1895 5919 5765 5856 2 1 5859 QDFFRBN $T=1037880 819960 0 180 $X=1026100 $Y=814540
X1896 5942 5765 5805 2 1 5882 QDFFRBN $T=1042220 799800 1 180 $X=1030440 $Y=799420
X1897 5893 1150 5853 2 1 5931 QDFFRBN $T=1031060 749400 0 0 $X=1031060 $Y=749020
X1898 5901 5765 5564 2 1 5921 QDFFRBN $T=1033540 840120 0 0 $X=1033540 $Y=839740
X1899 5912 5765 5564 2 1 5966 QDFFRBN $T=1034160 830040 1 0 $X=1034160 $Y=824620
X1900 5913 1146 1183 2 1 5920 QDFFRBN $T=1034160 870360 0 0 $X=1034160 $Y=869980
X1901 5918 5765 5949 2 1 5933 QDFFRBN $T=1034780 789720 0 0 $X=1034780 $Y=789340
X1902 5932 1150 5819 2 1 5897 QDFFRBN $T=1048420 759480 1 180 $X=1036640 $Y=759100
X1903 5883 1146 1183 2 1 5914 QDFFRBN $T=1037260 880440 0 0 $X=1037260 $Y=880060
X1904 5905 1146 1179 2 1 1167 QDFFRBN $T=1049040 900600 0 180 $X=1037260 $Y=895180
X1905 5989 5765 5949 2 1 5936 QDFFRBN $T=1049660 789720 0 180 $X=1037880 $Y=784300
X1906 5938 1146 1183 2 1 5929 QDFFRBN $T=1037880 890520 0 0 $X=1037880 $Y=890140
X1907 6010 5765 5943 2 1 5960 QDFFRBN $T=1054620 799800 0 180 $X=1042840 $Y=794380
X1908 6031 1150 1180 2 1 5973 QDFFRBN $T=1057100 729240 0 180 $X=1045320 $Y=723820
X1909 6013 5765 5949 2 1 5975 QDFFRBN $T=1057100 769560 1 180 $X=1045320 $Y=769180
X1910 6027 5765 5943 2 1 5979 QDFFRBN $T=1057720 840120 1 180 $X=1045940 $Y=839740
X1911 5983 1150 1180 2 1 5911 QDFFRBN $T=1058340 729240 1 180 $X=1046560 $Y=728860
X1912 6038 1146 6004 2 1 5984 QDFFRBN $T=1058960 850200 0 180 $X=1047180 $Y=844780
X1913 6049 1150 5974 2 1 5986 QDFFRBN $T=1059580 749400 1 180 $X=1047800 $Y=749020
X1914 5985 1146 6017 2 1 5957 QDFFRBN $T=1049660 860280 0 0 $X=1049660 $Y=859900
X1915 6007 1146 1183 2 1 6008 QDFFRBN $T=1050900 900600 1 0 $X=1050900 $Y=895180
X1916 6019 5765 5949 2 1 6006 QDFFRBN $T=1063300 769560 0 180 $X=1051520 $Y=764140
X1917 6009 5765 6033 2 1 6028 QDFFRBN $T=1052140 789720 1 0 $X=1052140 $Y=784300
X1918 6066 5765 6033 2 1 6011 QDFFRBN $T=1064540 799800 1 180 $X=1052760 $Y=799420
X1919 6021 5765 6003 2 1 5990 QDFFRBN $T=1054000 819960 1 0 $X=1054000 $Y=814540
X1920 6034 5765 6004 2 1 6037 QDFFRBN $T=1055860 830040 0 0 $X=1055860 $Y=829660
X1921 6035 5765 6033 2 1 6056 QDFFRBN $T=1056480 799800 1 0 $X=1056480 $Y=794380
X1922 6043 5765 6003 2 1 6062 QDFFRBN $T=1057720 840120 0 0 $X=1057720 $Y=839740
X1923 6044 1146 6017 2 1 6094 QDFFRBN $T=1057720 880440 0 0 $X=1057720 $Y=880060
X1924 6106 1146 6017 2 1 6055 QDFFRBN $T=1071980 890520 0 180 $X=1060200 $Y=885100
X1925 6059 1146 6017 2 1 6015 QDFFRBN $T=1060820 870360 1 0 $X=1060820 $Y=864940
X1926 6097 5765 5974 2 1 6067 QDFFRBN $T=1075080 759480 1 180 $X=1063300 $Y=759100
X1927 6074 1150 5974 2 1 1197 QDFFRBN $T=1063920 739320 1 0 $X=1063920 $Y=733900
X1928 6112 5765 6088 2 1 6075 QDFFRBN $T=1076320 769560 0 180 $X=1064540 $Y=764140
X1929 6083 1146 6128 2 1 6135 QDFFRBN $T=1066400 860280 0 0 $X=1066400 $Y=859900
X1930 6087 5765 6123 2 1 6103 QDFFRBN $T=1067020 799800 0 0 $X=1067020 $Y=799420
X1931 6132 5765 6033 2 1 6054 QDFFRBN $T=1079420 779640 1 180 $X=1067640 $Y=779260
X1932 6137 1150 5974 2 1 6090 QDFFRBN $T=1080040 739320 1 180 $X=1068260 $Y=738940
X1933 6141 5765 6088 2 1 6092 QDFFRBN $T=1080040 769560 1 180 $X=1068260 $Y=769180
X1934 6101 1146 6127 2 1 6133 QDFFRBN $T=1069500 840120 0 0 $X=1069500 $Y=839740
X1935 6111 1146 1216 2 1 1222 QDFFRBN $T=1070740 880440 0 0 $X=1070740 $Y=880060
X1936 6114 1150 6146 2 1 6120 QDFFRBN $T=1071360 749400 1 0 $X=1071360 $Y=743980
X1937 6115 5765 6127 2 1 6085 QDFFRBN $T=1071360 830040 0 0 $X=1071360 $Y=829660
X1938 6117 5765 6123 2 1 6125 QDFFRBN $T=1072600 819960 1 0 $X=1072600 $Y=814540
X1939 6167 1146 6017 2 1 1207 QDFFRBN $T=1086860 890520 0 180 $X=1075080 $Y=885100
X1940 6152 1150 6146 2 1 1214 QDFFRBN $T=1091820 739320 0 180 $X=1080040 $Y=733900
X1941 6198 1146 6128 2 1 6156 QDFFRBN $T=1092440 860280 1 180 $X=1080660 $Y=859900
X1942 6159 1146 1216 2 1 1225 QDFFRBN $T=1080660 900600 1 0 $X=1080660 $Y=895180
X1943 6208 5765 6123 2 1 6160 QDFFRBN $T=1093060 809880 1 180 $X=1081280 $Y=809500
X1944 6213 1150 6146 2 1 1221 QDFFRBN $T=1093680 729240 1 180 $X=1081900 $Y=728860
X1945 6214 1150 6146 2 1 6163 QDFFRBN $T=1093680 739320 1 180 $X=1081900 $Y=738940
X1946 6212 5765 6088 2 1 6157 QDFFRBN $T=1093680 769560 1 180 $X=1081900 $Y=769180
X1947 6166 1146 6206 2 1 6185 QDFFRBN $T=1083140 880440 0 0 $X=1083140 $Y=880060
X1948 6219 5765 6140 2 1 6174 QDFFRBN $T=1096780 779640 1 180 $X=1085000 $Y=779260
X1949 6182 5765 6188 2 1 6205 QDFFRBN $T=1085620 819960 1 0 $X=1085620 $Y=814540
X1950 6237 5765 6210 2 1 6196 QDFFRBN $T=1100500 799800 0 180 $X=1088720 $Y=794380
X1951 6200 5765 6188 2 1 6204 QDFFRBN $T=1089340 819960 0 0 $X=1089340 $Y=819580
X1952 6257 1146 6206 2 1 6193 QDFFRBN $T=1101740 890520 0 180 $X=1089960 $Y=885100
X1953 6215 5765 6128 2 1 6238 QDFFRBN $T=1091820 840120 0 0 $X=1091820 $Y=839740
X1954 6271 1146 6206 2 1 1228 QDFFRBN $T=1104840 890520 1 180 $X=1093060 $Y=890140
X1955 6279 1150 6224 2 1 6225 QDFFRBN $T=1106080 739320 1 180 $X=1094300 $Y=738940
X1956 6241 1146 6128 2 1 6207 QDFFRBN $T=1106080 850200 0 180 $X=1094300 $Y=844780
X1957 6245 1146 6128 2 1 6211 QDFFRBN $T=1106080 870360 0 180 $X=1094300 $Y=864940
X1958 6230 1150 6224 2 1 6259 QDFFRBN $T=1094920 729240 0 0 $X=1094920 $Y=728860
X1959 6283 1150 6224 2 1 6227 QDFFRBN $T=1106700 749400 0 180 $X=1094920 $Y=743980
X1960 6274 5765 6210 2 1 6228 QDFFRBN $T=1106700 809880 1 180 $X=1094920 $Y=809500
X1961 6291 5765 6224 2 1 6232 QDFFRBN $T=1107320 769560 1 180 $X=1095540 $Y=769180
X1962 6294 5765 6224 2 1 6249 QDFFRBN $T=1110420 769560 0 180 $X=1098640 $Y=764140
X1963 6314 5765 6140 2 1 6250 QDFFRBN $T=1110420 779640 1 180 $X=1098640 $Y=779260
X1964 6264 1146 6251 2 1 6256 QDFFRBN $T=1100500 860280 1 0 $X=1100500 $Y=854860
X1965 6278 5765 6188 2 1 6254 QDFFRBN $T=1114140 799800 0 180 $X=1102360 $Y=794380
X1966 6288 5765 6251 2 1 6246 QDFFRBN $T=1114760 819960 1 180 $X=1102980 $Y=819580
X1967 6276 1146 1247 2 1 6324 QDFFRBN $T=1103600 900600 1 0 $X=1103600 $Y=895180
X1968 6346 5765 6210 2 1 6297 QDFFRBN $T=1118480 819960 0 180 $X=1106700 $Y=814540
X1969 6321 1146 6251 2 1 6263 QDFFRBN $T=1119100 850200 0 180 $X=1107320 $Y=844780
X1970 6327 1146 6206 2 1 6267 QDFFRBN $T=1125920 840120 1 180 $X=1114140 $Y=839740
X1971 6332 1150 6369 2 1 6310 QDFFRBN $T=1128400 739320 1 180 $X=1116620 $Y=738940
X1972 6366 5765 6210 2 1 6340 QDFFRBN $T=1128400 809880 1 180 $X=1116620 $Y=809500
X1973 6349 5765 6362 2 1 6290 QDFFRBN $T=1128400 830040 0 180 $X=1116620 $Y=824620
X1974 6350 1146 6251 2 1 6299 QDFFRBN $T=1128400 860280 0 180 $X=1116620 $Y=854860
X1975 6363 1146 1247 2 1 6323 QDFFRBN $T=1128400 880440 0 180 $X=1116620 $Y=875020
X1976 6364 1146 1247 2 1 1246 QDFFRBN $T=1128400 890520 1 180 $X=1116620 $Y=890140
X1977 6372 1146 1247 2 1 6316 QDFFRBN $T=1128400 900600 0 180 $X=1116620 $Y=895180
X1978 6368 1150 1253 2 1 6339 QDFFRBN $T=1129020 729240 1 180 $X=1117240 $Y=728860
X1979 6355 1150 6369 2 1 6319 QDFFRBN $T=1129020 749400 1 180 $X=1117240 $Y=749020
X1980 6356 5765 6369 2 1 6261 QDFFRBN $T=1129020 759480 1 180 $X=1117240 $Y=759100
X1981 6357 5765 6369 2 1 6313 QDFFRBN $T=1129020 769560 0 180 $X=1117240 $Y=764140
X1982 6348 5765 6140 2 1 6315 QDFFRBN $T=1129020 779640 1 180 $X=1117240 $Y=779260
X1983 6358 5765 6140 2 1 6220 QDFFRBN $T=1129020 789720 0 180 $X=1117240 $Y=784300
X1984 6365 5765 6210 2 1 6307 QDFFRBN $T=1129020 799800 0 180 $X=1117240 $Y=794380
X1985 6337 5765 6210 2 1 6302 QDFFRBN $T=1129020 799800 1 180 $X=1117240 $Y=799420
X1986 6318 5765 6251 2 1 6269 QDFFRBN $T=1129020 819960 1 180 $X=1117240 $Y=819580
X1987 6359 5765 6362 2 1 6296 QDFFRBN $T=1129020 830040 1 180 $X=1117240 $Y=829660
X1988 6373 1146 6362 2 1 6328 QDFFRBN $T=1129020 850200 1 180 $X=1117240 $Y=849820
X1989 6360 1146 6362 2 1 1245 QDFFRBN $T=1129020 870360 0 180 $X=1117240 $Y=864940
X1990 6361 1146 6362 2 1 6329 QDFFRBN $T=1129020 870360 1 180 $X=1117240 $Y=869980
X1991 6347 5765 6369 2 1 6317 QDFFRBN $T=1129640 769560 1 180 $X=1117860 $Y=769180
X1992 2398 1 2 2423 2427 2467 1306 ICV_4 $T=397420 830040 0 0 $X=397420 $Y=829660
X1993 312 1 2 321 2598 2618 1306 ICV_4 $T=427180 799800 1 0 $X=427180 $Y=794380
X1994 2601 1 2 2621 2627 2650 1306 ICV_4 $T=432760 819960 0 0 $X=432760 $Y=819580
X1995 2602 1 2 2622 2628 2651 1306 ICV_4 $T=432760 840120 1 0 $X=432760 $Y=834700
X1996 2669 1 2 2679 2709 2735 1306 ICV_4 $T=446400 840120 0 0 $X=446400 $Y=839740
X1997 341 1 2 350 352 357 1306 ICV_4 $T=447640 900600 1 0 $X=447640 $Y=895180
X1998 2727 1 2 2747 2751 2775 1306 ICV_4 $T=455700 759480 0 0 $X=455700 $Y=759100
X1999 2724 1 2 2749 2744 2755 1306 ICV_4 $T=458180 830040 1 0 $X=458180 $Y=824620
X2000 2676 1 2 2691 2741 373 1306 ICV_4 $T=459420 890520 0 0 $X=459420 $Y=890140
X2001 2759 1 2 2760 2789 2793 1306 ICV_4 $T=462520 769560 1 0 $X=462520 $Y=764140
X2002 2716 1 2 2776 2720 2719 1306 ICV_4 $T=465000 860280 0 0 $X=465000 $Y=859900
X2003 2778 1 2 2790 2740 2695 1306 ICV_4 $T=468100 890520 1 0 $X=468100 $Y=885100
X2004 2804 1 2 2812 2835 2836 1306 ICV_4 $T=471200 830040 1 0 $X=471200 $Y=824620
X2005 2806 1 2 2830 2884 2891 1306 ICV_4 $T=483600 779640 1 0 $X=483600 $Y=774220
X2006 390 1 2 2888 2908 2887 1306 ICV_4 $T=487320 890520 1 0 $X=487320 $Y=885100
X2007 2859 1 2 2872 2746 2837 1306 ICV_4 $T=489180 850200 0 0 $X=489180 $Y=849820
X2008 2880 1 2 2893 2889 2906 1306 ICV_4 $T=491660 850200 1 0 $X=491660 $Y=844780
X2009 2886 1 2 2926 2897 2959 1306 ICV_4 $T=494140 880440 0 0 $X=494140 $Y=880060
X2010 2979 1 2 2964 3027 2998 1306 ICV_4 $T=507160 789720 0 0 $X=507160 $Y=789340
X2011 3042 1 2 3064 3075 3098 1306 ICV_4 $T=515840 739320 1 0 $X=515840 $Y=733900
X2012 3056 1 2 3052 3065 3091 1306 ICV_4 $T=519560 779640 0 0 $X=519560 $Y=779260
X2013 3076 1 2 3070 3071 3106 1306 ICV_4 $T=523280 739320 0 0 $X=523280 $Y=738940
X2014 3122 1 2 3152 3145 3156 1306 ICV_4 $T=530100 799800 0 0 $X=530100 $Y=799420
X2015 3139 1 2 3185 3147 3153 1306 ICV_4 $T=540640 840120 0 0 $X=540640 $Y=839740
X2016 3218 1 2 3245 3249 3267 1306 ICV_4 $T=549320 870360 1 0 $X=549320 $Y=864940
X2017 3219 1 2 3220 3154 3144 1306 ICV_4 $T=549940 759480 0 0 $X=549940 $Y=759100
X2018 3264 1 2 3265 3292 3320 1306 ICV_4 $T=558620 789720 0 0 $X=558620 $Y=789340
X2019 3266 1 2 3217 3222 3244 1306 ICV_4 $T=558620 830040 0 0 $X=558620 $Y=829660
X2020 3353 1 2 3347 3386 3360 1306 ICV_4 $T=573500 860280 0 0 $X=573500 $Y=859900
X2021 492 1 2 3323 3409 3380 1306 ICV_4 $T=575980 890520 1 0 $X=575980 $Y=885100
X2022 3423 1 2 3442 536 3445 1306 ICV_4 $T=586520 890520 0 0 $X=586520 $Y=890140
X2023 3399 1 2 3426 3449 3459 1306 ICV_4 $T=593340 819960 1 0 $X=593340 $Y=814540
X2024 3465 1 2 3474 3489 3530 1306 ICV_4 $T=600780 850200 1 0 $X=600780 $Y=844780
X2025 3525 1 2 3543 3521 3545 1306 ICV_4 $T=604500 880440 1 0 $X=604500 $Y=875020
X2026 3497 1 2 3534 3552 3571 1306 ICV_4 $T=606360 819960 1 0 $X=606360 $Y=814540
X2027 3610 1 2 3640 592 598 1306 ICV_4 $T=623720 729240 1 0 $X=623720 $Y=723820
X2028 3602 1 2 3642 3634 3665 1306 ICV_4 $T=624340 759480 0 0 $X=624340 $Y=759100
X2029 587 1 2 3660 3661 3684 1306 ICV_4 $T=627440 890520 0 0 $X=627440 $Y=890140
X2030 3675 1 2 3696 3701 3720 1306 ICV_4 $T=636120 850200 1 0 $X=636120 $Y=844780
X2031 3682 1 2 3699 3670 3704 1306 ICV_4 $T=636740 759480 0 0 $X=636740 $Y=759100
X2032 3709 1 2 3719 3695 3759 1306 ICV_4 $T=642940 789720 1 0 $X=642940 $Y=784300
X2033 3728 1 2 3743 3751 3744 1306 ICV_4 $T=646660 860280 1 0 $X=646660 $Y=854860
X2034 3754 1 2 3749 3780 3806 1306 ICV_4 $T=652240 769560 0 0 $X=652240 $Y=769180
X2035 3790 1 2 3815 3819 3818 1306 ICV_4 $T=659680 759480 0 0 $X=659680 $Y=759100
X2036 3758 1 2 3738 3812 3807 1306 ICV_4 $T=662780 840120 1 0 $X=662780 $Y=834700
X2037 3865 1 2 3809 3861 3850 1306 ICV_4 $T=673940 819960 0 0 $X=673940 $Y=819580
X2038 683 1 2 3874 684 3901 1306 ICV_4 $T=676420 880440 0 0 $X=676420 $Y=880060
X2039 3826 1 2 3835 3929 3970 1306 ICV_4 $T=684480 779640 0 0 $X=684480 $Y=779260
X2040 3961 1 2 3939 3977 4001 1306 ICV_4 $T=693780 789720 1 0 $X=693780 $Y=784300
X2041 3932 1 2 3962 4056 4049 1306 ICV_4 $T=701220 870360 1 0 $X=701220 $Y=864940
X2042 3949 1 2 3992 3860 3948 1306 ICV_4 $T=706180 779640 0 0 $X=706180 $Y=779260
X2043 4082 1 2 4084 4077 4074 1306 ICV_4 $T=730980 809880 0 0 $X=730980 $Y=809500
X2044 4258 1 2 4281 4200 4306 1306 ICV_4 $T=744000 840120 0 0 $X=744000 $Y=839740
X2045 4247 1 2 4257 824 831 1306 ICV_4 $T=745240 890520 0 0 $X=745240 $Y=890140
X2046 4313 1 2 4336 4341 4363 1306 ICV_4 $T=755780 870360 1 0 $X=755780 $Y=864940
X2047 4335 1 2 4356 4358 4371 1306 ICV_4 $T=759500 789720 1 0 $X=759500 $Y=784300
X2048 4401 1 2 4404 4390 4411 1306 ICV_4 $T=771900 830040 1 0 $X=771900 $Y=824620
X2049 863 1 2 872 4452 4466 1306 ICV_4 $T=773140 900600 1 0 $X=773140 $Y=895180
X2050 4472 1 2 4502 4504 4507 1306 ICV_4 $T=783680 779640 1 0 $X=783680 $Y=774220
X2051 4501 1 2 4528 900 905 1306 ICV_4 $T=788020 739320 1 0 $X=788020 $Y=733900
X2052 4522 1 2 4548 4554 4579 1306 ICV_4 $T=791120 819960 1 0 $X=791120 $Y=814540
X2053 4531 1 2 4563 4567 4599 1306 ICV_4 $T=792980 819960 0 0 $X=792980 $Y=819580
X2054 4565 1 2 4594 4598 4625 1306 ICV_4 $T=797940 799800 0 0 $X=797940 $Y=799420
X2055 4597 1 2 4622 4616 4632 1306 ICV_4 $T=802900 759480 0 0 $X=802900 $Y=759100
X2056 4601 1 2 4647 942 950 1306 ICV_4 $T=816540 880440 0 0 $X=816540 $Y=880060
X2057 4691 1 2 4724 4723 4747 1306 ICV_4 $T=819640 729240 0 0 $X=819640 $Y=728860
X2058 4735 1 2 4762 4761 4794 1306 ICV_4 $T=825840 840120 0 0 $X=825840 $Y=839740
X2059 953 1 2 955 958 962 1306 ICV_4 $T=830180 880440 0 0 $X=830180 $Y=880060
X2060 4817 1 2 4827 4818 4834 1306 ICV_4 $T=840720 729240 1 0 $X=840720 $Y=723820
X2061 4808 1 2 4829 4848 4841 1306 ICV_4 $T=841340 769560 0 0 $X=841340 $Y=769180
X2062 4875 1 2 4904 4906 4925 1306 ICV_4 $T=851260 769560 0 0 $X=851260 $Y=769180
X2063 4898 1 2 4920 4922 4923 1306 ICV_4 $T=854980 729240 1 0 $X=854980 $Y=723820
X2064 4942 1 2 4939 4969 4997 1306 ICV_4 $T=864280 860280 1 0 $X=864280 $Y=854860
X2065 4943 1 2 4935 4980 4995 1306 ICV_4 $T=866760 799800 1 0 $X=866760 $Y=794380
X2066 4805 1 2 4828 4956 4998 1306 ICV_4 $T=868620 830040 1 0 $X=868620 $Y=824620
X2067 4973 1 2 4999 997 5029 1306 ICV_4 $T=869860 900600 1 0 $X=869860 $Y=895180
X2068 5023 1 2 5027 5060 5066 1306 ICV_4 $T=879780 789720 1 0 $X=879780 $Y=784300
X2069 4926 1 2 4909 5069 5079 1306 ICV_4 $T=882880 749400 1 0 $X=882880 $Y=743980
X2070 5065 1 2 5072 5047 5090 1306 ICV_4 $T=885360 860280 1 0 $X=885360 $Y=854860
X2071 5149 1 2 5148 5137 5152 1306 ICV_4 $T=900860 739320 0 0 $X=900860 $Y=738940
X2072 5084 1 2 5118 5157 5190 1306 ICV_4 $T=905200 860280 0 0 $X=905200 $Y=859900
X2073 5153 1 2 5163 5166 5173 1306 ICV_4 $T=908920 769560 1 0 $X=908920 $Y=764140
X2074 5203 1 2 5204 5193 5220 1306 ICV_4 $T=910780 819960 1 0 $X=910780 $Y=814540
X2075 5255 1 2 5273 5265 5278 1306 ICV_4 $T=923180 729240 0 0 $X=923180 $Y=728860
X2076 5264 1 2 5298 5305 5313 1306 ICV_4 $T=926280 890520 1 0 $X=926280 $Y=885100
X2077 5237 1 2 5352 5358 5365 1306 ICV_4 $T=934340 779640 1 0 $X=934340 $Y=774220
X2078 5301 1 2 5322 5299 5290 1306 ICV_4 $T=934960 819960 1 0 $X=934960 $Y=814540
X2079 5371 1 2 5357 5405 5344 1306 ICV_4 $T=942400 739320 1 0 $X=942400 $Y=733900
X2080 5310 1 2 5339 5377 5281 1306 ICV_4 $T=943640 769560 0 0 $X=943640 $Y=769180
X2081 5442 1 2 5447 5474 5493 1306 ICV_4 $T=956660 739320 0 0 $X=956660 $Y=738940
X2082 5547 1 2 5546 5573 5556 1306 ICV_4 $T=970300 870360 1 0 $X=970300 $Y=864940
X2083 5599 1 2 5609 5603 5610 1306 ICV_4 $T=983320 819960 0 0 $X=983320 $Y=819580
X2084 5579 1 2 5597 5658 5668 1306 ICV_4 $T=992620 870360 1 0 $X=992620 $Y=864940
X2085 5692 1 2 5731 5682 5740 1306 ICV_4 $T=999440 769560 0 0 $X=999440 $Y=769180
X2086 5532 1 2 5576 5673 5654 1306 ICV_4 $T=1001300 749400 0 0 $X=1001300 $Y=749020
X2087 5401 1 2 5441 5540 5613 1306 ICV_4 $T=1018660 870360 0 0 $X=1018660 $Y=869980
X2088 5859 1 2 5892 5921 5922 1306 ICV_4 $T=1031060 840120 1 0 $X=1031060 $Y=834700
X2089 5046 1 2 5074 1175 1181 1306 ICV_4 $T=1032300 870360 1 0 $X=1032300 $Y=864940
X2090 5854 1 2 5823 5882 5927 1306 ICV_4 $T=1033540 809880 1 0 $X=1033540 $Y=804460
X2091 5979 1 2 5997 6015 6042 1306 ICV_4 $T=1048420 870360 0 0 $X=1048420 $Y=869980
X2092 5975 1 2 6001 6028 6051 1306 ICV_4 $T=1050280 779640 1 0 $X=1050280 $Y=774220
X2093 5641 1 2 5669 4936 4996 1306 ICV_4 $T=1058340 840120 1 0 $X=1058340 $Y=834700
X2094 6125 1 2 6143 6129 6154 1306 ICV_4 $T=1074460 789720 0 0 $X=1074460 $Y=789340
X2095 6135 1 2 6144 6156 6173 1306 ICV_4 $T=1076940 870360 0 0 $X=1076940 $Y=869980
X2096 6163 1 2 6191 6186 6195 1306 ICV_4 $T=1083760 749400 1 0 $X=1083760 $Y=743980
X2097 6196 1 2 6217 6160 6240 1306 ICV_4 $T=1092440 789720 1 0 $X=1092440 $Y=784300
X2098 6220 1 2 6244 1234 1237 1306 ICV_4 $T=1093060 739320 1 0 $X=1093060 $Y=733900
X2099 6207 1 2 6221 6211 6222 1306 ICV_4 $T=1093060 870360 0 0 $X=1093060 $Y=869980
X2100 6238 1 2 6252 6246 6266 1306 ICV_4 $T=1096780 830040 0 0 $X=1096780 $Y=829660
X2101 6157 1 2 6236 6249 6270 1306 ICV_4 $T=1097400 759480 0 0 $X=1097400 $Y=759100
X2102 6232 1 2 6272 6254 6262 1306 ICV_4 $T=1102980 789720 1 0 $X=1102980 $Y=784300
X2103 6171 1 2 6197 6204 6233 1306 ICV_4 $T=1106700 830040 0 0 $X=1106700 $Y=829660
X2104 6250 1 2 6277 6307 6342 1306 ICV_4 $T=1114140 789720 0 0 $X=1114140 $Y=789340
X2105 6310 1 2 6353 6322 6333 1306 ICV_4 $T=1116620 739320 1 0 $X=1116620 $Y=733900
X2106 6313 1 2 6336 6261 6335 1306 ICV_4 $T=1116620 759480 1 0 $X=1116620 $Y=754060
X2107 6296 1 2 6331 6290 6320 1306 ICV_4 $T=1116620 840120 1 0 $X=1116620 $Y=834700
X2108 6263 1 2 6300 6329 6338 1306 ICV_4 $T=1116620 860280 0 0 $X=1116620 $Y=859900
X2109 6324 1 2 6344 1254 1255 1306 ICV_4 $T=1116620 890520 1 0 $X=1116620 $Y=885100
X2110 6297 1 2 6309 6340 6343 1306 ICV_4 $T=1117240 809880 1 0 $X=1117240 $Y=804460
X2111 6339 1 2 6345 1050 5351 1306 ICV_4 $T=1118480 729240 1 0 $X=1118480 $Y=723820
X2112 6315 1 2 6326 6174 6175 1306 ICV_4 $T=1118480 779640 1 0 $X=1118480 $Y=774220
X2113 6205 1 2 6203 6267 6303 1306 ICV_4 $T=1118480 819960 1 0 $X=1118480 $Y=814540
X2114 99 1655 2 1 1588 90 MUX2 $T=287060 729240 0 180 $X=282720 $Y=723820
X2115 2001 2044 2 1 204 1690 MUX2 $T=346580 799800 1 0 $X=346580 $Y=794380
X2116 1993 2067 2 1 2098 1955 MUX2 $T=347200 789720 0 0 $X=347200 $Y=789340
X2117 198 2044 2 1 2155 177 MUX2 $T=355260 799800 0 0 $X=355260 $Y=799420
X2118 215 2044 2 1 2186 218 MUX2 $T=361460 799800 1 0 $X=361460 $Y=794380
X2119 241 2194 2 1 2281 1969 MUX2 $T=376340 799800 1 0 $X=376340 $Y=794380
X2120 242 2194 2 1 2293 2260 MUX2 $T=377580 789720 1 0 $X=377580 $Y=784300
X2121 2648 2656 2 1 2585 2630 MUX2 $T=442680 799800 0 180 $X=438340 $Y=794380
X2122 2574 331 2 1 2664 2652 MUX2 $T=440200 880440 0 0 $X=440200 $Y=880060
X2123 340 331 2 1 329 336 MUX2 $T=445160 900600 0 180 $X=440820 $Y=895180
X2124 2644 2656 2 1 2590 2155 MUX2 $T=446400 789720 0 180 $X=442060 $Y=784300
X2125 2579 2670 2 1 2600 2649 MUX2 $T=446400 809880 1 180 $X=442060 $Y=809500
X2126 2671 2692 2 1 2593 2155 MUX2 $T=447020 779640 1 180 $X=442680 $Y=779260
X2127 2679 2678 2 1 2611 338 MUX2 $T=447020 840120 0 180 $X=442680 $Y=834700
X2128 2509 2684 2 1 2623 2652 MUX2 $T=447020 870360 0 180 $X=442680 $Y=864940
X2129 2687 2692 2 1 2661 2660 MUX2 $T=448880 779640 0 180 $X=444540 $Y=774220
X2130 2617 2670 2 1 2591 2155 MUX2 $T=448880 809880 0 180 $X=444540 $Y=804460
X2131 2691 344 2 1 2604 2652 MUX2 $T=448880 890520 0 180 $X=444540 $Y=885100
X2132 2467 2680 2 1 2594 2649 MUX2 $T=452600 840120 0 180 $X=448260 $Y=834700
X2133 2622 2678 2 1 2613 2649 MUX2 $T=452600 850200 0 180 $X=448260 $Y=844780
X2134 2618 2656 2 1 2675 2712 MUX2 $T=448880 799800 1 0 $X=448880 $Y=794380
X2135 2695 331 2 1 2685 345 MUX2 $T=448880 890520 1 0 $X=448880 $Y=885100
X2136 2527 2680 2 1 2730 349 MUX2 $T=450120 830040 0 0 $X=450120 $Y=829660
X2137 2719 2717 2 1 2657 345 MUX2 $T=455080 870360 0 180 $X=450740 $Y=864940
X2138 2731 2692 2 1 2707 2712 MUX2 $T=456940 779640 1 180 $X=452600 $Y=779260
X2139 2735 2678 2 1 2681 349 MUX2 $T=458180 850200 0 180 $X=453840 $Y=844780
X2140 2749 2670 2 1 2696 349 MUX2 $T=458800 809880 0 180 $X=454460 $Y=804460
X2141 2760 2656 2 1 2723 2706 MUX2 $T=463140 779640 1 180 $X=458800 $Y=779260
X2142 2651 2678 2 1 2766 2706 MUX2 $T=458800 850200 1 0 $X=458800 $Y=844780
X2143 2776 2773 2 1 2748 345 MUX2 $T=464380 860280 0 180 $X=460040 $Y=854860
X2144 2755 2670 2 1 2777 2706 MUX2 $T=461900 809880 1 0 $X=461900 $Y=804460
X2145 2793 2692 2 1 2738 2706 MUX2 $T=468100 779640 0 180 $X=463760 $Y=774220
X2146 2800 2678 2 1 2768 365 MUX2 $T=468100 850200 0 180 $X=463760 $Y=844780
X2147 2588 2680 2 1 2753 2706 MUX2 $T=468720 830040 1 180 $X=464380 $Y=829660
X2148 2650 2670 2 1 2767 365 MUX2 $T=471820 809880 0 180 $X=467480 $Y=804460
X2149 2812 2680 2 1 2734 365 MUX2 $T=471820 840120 0 180 $X=467480 $Y=834700
X2150 2790 368 2 1 2813 2816 MUX2 $T=467480 880440 0 0 $X=467480 $Y=880060
X2151 2815 368 2 1 2791 370 MUX2 $T=472440 870360 1 180 $X=468100 $Y=869980
X2152 2558 2656 2 1 2825 2794 MUX2 $T=470580 779640 0 0 $X=470580 $Y=779260
X2153 2832 2678 2 1 2802 370 MUX2 $T=475540 840120 1 180 $X=471200 $Y=839740
X2154 2836 2680 2 1 2772 2299 MUX2 $T=476160 830040 1 180 $X=471820 $Y=829660
X2155 2705 2841 2 1 2826 2299 MUX2 $T=478640 809880 0 180 $X=474300 $Y=804460
X2156 2830 2692 2 1 2854 2794 MUX2 $T=474920 779640 0 0 $X=474920 $Y=779260
X2157 2848 380 2 1 2823 378 MUX2 $T=479260 900600 0 180 $X=474920 $Y=895180
X2158 2837 380 2 1 2851 2652 MUX2 $T=475540 880440 0 0 $X=475540 $Y=880060
X2159 2846 2867 2 1 2803 2794 MUX2 $T=482980 759480 1 180 $X=478640 $Y=759100
X2160 2872 2717 2 1 2788 2852 MUX2 $T=484220 860280 1 180 $X=479880 $Y=859900
X2161 2883 2867 2 1 2809 2660 MUX2 $T=486700 749400 0 180 $X=482360 $Y=743980
X2162 2737 2867 2 1 2810 2898 MUX2 $T=482360 749400 0 0 $X=482360 $Y=749020
X2163 2863 2845 2 1 2878 2871 MUX2 $T=482360 830040 0 0 $X=482360 $Y=829660
X2164 2887 394 2 1 2870 370 MUX2 $T=487940 880440 1 180 $X=483600 $Y=880060
X2165 2891 2841 2 1 2829 2871 MUX2 $T=488560 809880 1 180 $X=484220 $Y=809500
X2166 2875 2692 2 1 2865 2831 MUX2 $T=485460 769560 1 0 $X=485460 $Y=764140
X2167 2904 2876 2 1 2877 2160 MUX2 $T=491040 789720 0 180 $X=486700 $Y=784300
X2168 2906 2866 2 1 2862 2871 MUX2 $T=491040 830040 1 180 $X=486700 $Y=829660
X2169 2888 394 2 1 398 378 MUX2 $T=487320 900600 1 0 $X=487320 $Y=895180
X2170 2817 2867 2 1 2911 2155 MUX2 $T=487940 749400 1 0 $X=487940 $Y=743980
X2171 2925 2867 2 1 2868 2831 MUX2 $T=494760 749400 1 180 $X=490420 $Y=749020
X2172 405 2933 2 1 2864 401 MUX2 $T=498480 749400 0 180 $X=494140 $Y=743980
X2173 2939 2933 2 1 2873 402 MUX2 $T=498480 769560 0 180 $X=494140 $Y=764140
X2174 2921 2845 2 1 2942 2952 MUX2 $T=494760 830040 1 0 $X=494760 $Y=824620
X2175 2926 380 2 1 2938 2949 MUX2 $T=495380 870360 0 0 $X=495380 $Y=869980
X2176 2940 2876 2 1 2961 2963 MUX2 $T=497860 779640 0 0 $X=497860 $Y=779260
X2177 2964 2874 2 1 2909 2580 MUX2 $T=502820 799800 1 180 $X=498480 $Y=799420
X2178 2953 2933 2 1 413 409 MUX2 $T=499720 729240 1 0 $X=499720 $Y=723820
X2179 2982 2933 2 1 2958 2712 MUX2 $T=505300 769560 0 180 $X=500960 $Y=764140
X2180 2996 2867 2 1 2968 2242 MUX2 $T=507160 749400 1 180 $X=502820 $Y=749020
X2181 3000 2841 2 1 2962 2952 MUX2 $T=507780 809880 1 180 $X=503440 $Y=809500
X2182 418 2933 2 1 2935 428 MUX2 $T=508400 729240 1 0 $X=508400 $Y=723820
X2183 3052 2977 2 1 3002 3015 MUX2 $T=518320 789720 0 180 $X=513980 $Y=784300
X2184 3085 3074 2 1 3047 402 MUX2 $T=523900 769560 0 180 $X=519560 $Y=764140
X2185 3073 2882 2 1 3080 3094 MUX2 $T=520800 860280 1 0 $X=520800 $Y=854860
X2186 3106 3109 2 1 3012 402 MUX2 $T=525760 749400 1 180 $X=521420 $Y=749020
X2187 2275 3095 2 1 3063 2871 MUX2 $T=525760 850200 1 180 $X=521420 $Y=849820
X2188 3086 437 2 1 3107 3094 MUX2 $T=523280 880440 0 0 $X=523280 $Y=880060
X2189 3064 3109 2 1 3024 409 MUX2 $T=528860 729240 1 180 $X=524520 $Y=728860
X2190 3091 2977 2 1 3119 2234 MUX2 $T=524520 789720 1 0 $X=524520 $Y=784300
X2191 3123 2937 2 1 3079 2306 MUX2 $T=530100 799800 1 180 $X=525760 $Y=799420
X2192 3090 3093 2 1 3082 2580 MUX2 $T=525760 830040 0 0 $X=525760 $Y=829660
X2193 3125 2882 2 1 3097 3101 MUX2 $T=530100 850200 1 180 $X=525760 $Y=849820
X2194 3159 3109 2 1 3096 426 MUX2 $T=532580 749400 1 180 $X=528240 $Y=749020
X2195 3144 3074 2 1 3089 426 MUX2 $T=533200 759480 1 180 $X=528860 $Y=759100
X2196 3153 3093 2 1 3103 3101 MUX2 $T=534440 830040 1 180 $X=530100 $Y=829660
X2197 3134 3109 2 1 450 428 MUX2 $T=531960 729240 0 0 $X=531960 $Y=728860
X2198 448 3109 2 1 3179 401 MUX2 $T=536920 729240 1 0 $X=536920 $Y=723820
X2199 3183 3074 2 1 3200 459 MUX2 $T=540640 759480 0 0 $X=540640 $Y=759100
X2200 3185 3068 2 1 3201 3101 MUX2 $T=540640 850200 0 0 $X=540640 $Y=849820
X2201 3220 3061 2 1 3198 2963 MUX2 $T=550560 769560 1 180 $X=546220 $Y=769180
X2202 3117 3004 2 1 3221 2306 MUX2 $T=546220 799800 0 0 $X=546220 $Y=799420
X2203 465 3109 2 1 3239 459 MUX2 $T=549320 749400 0 0 $X=549320 $Y=749020
X2204 3217 3215 2 1 3241 2580 MUX2 $T=549320 830040 0 0 $X=549320 $Y=829660
X2205 3205 3190 2 1 3193 459 MUX2 $T=554900 779640 1 180 $X=550560 $Y=779260
X2206 3244 3247 2 1 3260 3094 MUX2 $T=553660 819960 0 0 $X=553660 $Y=819580
X2207 3265 3256 2 1 3243 2306 MUX2 $T=559240 799800 0 180 $X=554900 $Y=794380
X2208 3270 3271 2 1 3216 3253 MUX2 $T=559240 870360 1 180 $X=554900 $Y=869980
X2209 3275 3252 2 1 3236 474 MUX2 $T=560480 739320 0 180 $X=556140 $Y=733900
X2210 3245 466 2 1 3305 3186 MUX2 $T=556140 890520 1 0 $X=556140 $Y=885100
X2211 3282 3271 2 1 3191 3186 MUX2 $T=561100 880440 1 180 $X=556760 $Y=880060
X2212 3307 3204 2 1 3237 3233 MUX2 $T=566060 749400 1 180 $X=561720 $Y=749020
X2213 3267 466 2 1 3212 3318 MUX2 $T=562960 860280 1 0 $X=562960 $Y=854860
X2214 3299 3247 2 1 3238 3317 MUX2 $T=563580 840120 0 0 $X=563580 $Y=839740
X2215 3323 480 2 1 483 481 MUX2 $T=568540 890520 1 180 $X=564200 $Y=890140
X2216 3320 3190 2 1 3338 3343 MUX2 $T=567300 779640 0 0 $X=567300 $Y=779260
X2217 3339 3345 2 1 3359 3285 MUX2 $T=571020 819960 1 0 $X=571020 $Y=814540
X2218 3360 3345 2 1 3340 3318 MUX2 $T=575360 860280 0 180 $X=571020 $Y=854860
X2219 3347 3345 2 1 3376 3352 MUX2 $T=573500 850200 1 0 $X=573500 $Y=844780
X2220 3380 511 2 1 3354 3186 MUX2 $T=578460 880440 1 180 $X=574120 $Y=880060
X2221 3358 3256 2 1 3377 3384 MUX2 $T=574740 799800 1 0 $X=574740 $Y=794380
X2222 517 3413 2 1 3306 2234 MUX2 $T=582800 769560 0 180 $X=578460 $Y=764140
X2223 3400 3345 2 1 3390 3316 MUX2 $T=579700 840120 1 0 $X=579700 $Y=834700
X2224 2747 3432 2 1 3349 3318 MUX2 $T=589620 850200 1 180 $X=585280 $Y=849820
X2225 3445 538 2 1 543 481 MUX2 $T=591480 900600 1 0 $X=591480 $Y=895180
X2226 3446 3204 2 1 3466 3467 MUX2 $T=592100 769560 1 0 $X=592100 $Y=764140
X2227 542 3204 2 1 3478 3482 MUX2 $T=594580 749400 0 0 $X=594580 $Y=749020
X2228 3459 3464 2 1 3483 3285 MUX2 $T=594580 819960 0 0 $X=594580 $Y=819580
X2229 2551 538 2 1 3503 3186 MUX2 $T=598300 880440 0 0 $X=598300 $Y=880060
X2230 3452 3490 2 1 3518 3101 MUX2 $T=599540 769560 1 0 $X=599540 $Y=764140
X2231 3523 3527 2 1 3470 3101 MUX2 $T=605120 749400 1 180 $X=600780 $Y=749020
X2232 2775 3528 2 1 3508 3487 MUX2 $T=606360 789720 1 180 $X=602020 $Y=789340
X2233 553 554 2 1 3512 3511 MUX2 $T=606360 900600 0 180 $X=602020 $Y=895180
X2234 3534 3501 2 1 3514 3285 MUX2 $T=606980 819960 1 180 $X=602640 $Y=819580
X2235 3529 3549 2 1 3506 3487 MUX2 $T=610080 799800 1 180 $X=605740 $Y=799420
X2236 3551 3554 2 1 3515 545 MUX2 $T=611940 739320 1 180 $X=607600 $Y=738940
X2237 556 3490 2 1 3516 560 MUX2 $T=608840 779640 1 0 $X=608840 $Y=774220
X2238 3545 3485 2 1 3561 3566 MUX2 $T=609460 860280 0 0 $X=609460 $Y=859900
X2239 2570 3546 2 1 3578 3186 MUX2 $T=613180 880440 0 0 $X=613180 $Y=880060
X2240 3591 3563 2 1 3522 3562 MUX2 $T=619380 809880 0 180 $X=615040 $Y=804460
X2241 3442 3572 2 1 3616 3593 MUX2 $T=616900 880440 1 0 $X=616900 $Y=875020
X2242 3603 3584 2 1 3587 3562 MUX2 $T=622480 809880 1 180 $X=618140 $Y=809500
X2243 3447 563 2 1 576 3511 MUX2 $T=618140 900600 1 0 $X=618140 $Y=895180
X2244 3595 3572 2 1 3626 3566 MUX2 $T=620000 870360 1 0 $X=620000 $Y=864940
X2245 579 3484 2 1 3648 3652 MUX2 $T=625580 850200 0 0 $X=625580 $Y=849820
X2246 596 3655 2 1 3622 3482 MUX2 $T=631780 830040 1 180 $X=627440 $Y=829660
X2247 600 578 2 1 3649 3487 MUX2 $T=633640 769560 0 180 $X=629300 $Y=764140
X2248 3650 3647 2 1 3668 3562 MUX2 $T=629300 809880 0 0 $X=629300 $Y=809500
X2249 601 3669 2 1 3653 3566 MUX2 $T=634260 870360 0 180 $X=629920 $Y=864940
X2250 606 3679 2 1 3659 3467 MUX2 $T=636120 799800 0 180 $X=631780 $Y=794380
X2251 609 3647 2 1 3614 3482 MUX2 $T=636120 819960 1 180 $X=631780 $Y=819580
X2252 3571 3693 2 1 3604 3562 MUX2 $T=638600 819960 0 180 $X=634260 $Y=814540
X2253 3646 3655 2 1 3698 607 MUX2 $T=636120 860280 1 0 $X=636120 $Y=854860
X2254 619 3655 2 1 3671 3652 MUX2 $T=641700 840120 1 180 $X=637360 $Y=839740
X2255 3688 608 2 1 3702 3593 MUX2 $T=637360 880440 1 0 $X=637360 $Y=875020
X2256 3666 3647 2 1 3708 3652 MUX2 $T=637980 809880 0 0 $X=637980 $Y=809500
X2257 612 608 2 1 3711 3511 MUX2 $T=638600 900600 1 0 $X=638600 $Y=895180
X2258 3704 3554 2 1 3718 560 MUX2 $T=641700 749400 0 0 $X=641700 $Y=749020
X2259 3660 608 2 1 624 625 MUX2 $T=646660 890520 1 180 $X=642320 $Y=890140
X2260 3732 3706 2 1 3676 3713 MUX2 $T=647900 769560 1 180 $X=643560 $Y=769180
X2261 634 605 2 1 627 629 MUX2 $T=650380 729240 0 180 $X=646040 $Y=723820
X2262 3609 3724 2 1 3715 3738 MUX2 $T=646040 840120 1 0 $X=646040 $Y=834700
X2263 3684 637 2 1 3730 3511 MUX2 $T=651000 890520 1 180 $X=646660 $Y=890140
X2264 3744 3729 2 1 3710 3566 MUX2 $T=651620 870360 0 180 $X=647280 $Y=864940
X2265 640 637 2 1 633 625 MUX2 $T=651620 900600 0 180 $X=647280 $Y=895180
X2266 3749 3678 2 1 3733 3713 MUX2 $T=652240 769560 1 180 $X=647900 $Y=769180
X2267 3720 3655 2 1 3756 3764 MUX2 $T=648520 830040 0 0 $X=648520 $Y=829660
X2268 636 3606 2 1 3763 3713 MUX2 $T=651000 739320 0 0 $X=651000 $Y=738940
X2269 3759 3678 2 1 3741 3652 MUX2 $T=656580 779640 1 180 $X=652240 $Y=779260
X2270 3777 637 2 1 3752 3593 MUX2 $T=657200 880440 1 180 $X=652860 $Y=880060
X2271 3699 3693 2 1 3786 3713 MUX2 $T=655960 809880 0 0 $X=655960 $Y=809500
X2272 646 605 2 1 650 651 MUX2 $T=656580 729240 1 0 $X=656580 $Y=723820
X2273 3696 3737 2 1 3798 3764 MUX2 $T=656580 830040 0 0 $X=656580 $Y=829660
X2274 652 3606 2 1 3784 3692 MUX2 $T=662160 739320 1 180 $X=657820 $Y=738940
X2275 653 3679 2 1 3787 3713 MUX2 $T=662780 799800 0 180 $X=658440 $Y=794380
X2276 3818 3662 2 1 3799 402 MUX2 $T=665260 749400 0 180 $X=660920 $Y=743980
X2277 3801 3693 2 1 3760 3692 MUX2 $T=665880 789720 1 180 $X=661540 $Y=789340
X2278 3809 3808 2 1 3824 3609 MUX2 $T=662160 830040 0 0 $X=662160 $Y=829660
X2279 3830 3825 2 1 3804 3593 MUX2 $T=668360 880440 0 180 $X=664020 $Y=875020
X2280 668 3678 2 1 3820 3692 MUX2 $T=668980 769560 0 180 $X=664640 $Y=764140
X2281 3815 3662 2 1 3823 3692 MUX2 $T=669600 749400 0 180 $X=665260 $Y=743980
X2282 3581 3808 2 1 3788 3352 MUX2 $T=670220 850200 0 180 $X=665880 $Y=844780
X2283 3852 3678 2 1 3817 3829 MUX2 $T=671460 779640 0 180 $X=667120 $Y=774220
X2284 664 605 2 1 673 677 MUX2 $T=668360 729240 1 0 $X=668360 $Y=723820
X2285 3745 672 2 1 3805 3511 MUX2 $T=672700 890520 1 180 $X=668360 $Y=890140
X2286 674 3822 2 1 3768 651 MUX2 $T=673320 729240 1 180 $X=668980 $Y=728860
X2287 3835 3832 2 1 3855 3692 MUX2 $T=668980 789720 0 0 $X=668980 $Y=789340
X2288 3850 3828 2 1 3811 3829 MUX2 $T=673320 799800 1 180 $X=668980 $Y=799420
X2289 3834 672 2 1 3863 3318 MUX2 $T=670840 870360 1 0 $X=670840 $Y=864940
X2290 3879 3858 2 1 3843 3352 MUX2 $T=678280 850200 1 180 $X=673940 $Y=849820
X2291 3869 3706 2 1 3886 3829 MUX2 $T=675180 769560 0 0 $X=675180 $Y=769180
X2292 689 3822 2 1 3851 3875 MUX2 $T=681380 729240 1 180 $X=677040 $Y=728860
X2293 3743 3808 2 1 3882 3652 MUX2 $T=682620 840120 1 180 $X=678280 $Y=839740
X2294 3901 692 2 1 697 625 MUX2 $T=680760 900600 1 0 $X=680760 $Y=895180
X2295 3939 3832 2 1 3909 3910 MUX2 $T=688200 799800 0 180 $X=683860 $Y=794380
X2296 3923 3808 2 1 3938 654 MUX2 $T=685100 830040 0 0 $X=685100 $Y=829660
X2297 3924 3906 2 1 3945 3875 MUX2 $T=685720 749400 1 0 $X=685720 $Y=743980
X2298 3948 3947 2 1 3914 3910 MUX2 $T=690060 779640 0 180 $X=685720 $Y=774220
X2299 706 3956 2 1 3848 3593 MUX2 $T=691300 880440 0 180 $X=686960 $Y=875020
X2300 3975 3822 2 1 3927 3946 MUX2 $T=693780 729240 1 180 $X=689440 $Y=728860
X2301 711 3706 2 1 3908 3946 MUX2 $T=694400 779640 0 180 $X=690060 $Y=774220
X2302 3976 3828 2 1 3915 3910 MUX2 $T=694400 809880 0 180 $X=690060 $Y=804460
X2303 3992 3828 2 1 3883 3946 MUX2 $T=695640 789720 1 180 $X=691300 $Y=789340
X2304 3962 3956 2 1 3984 3318 MUX2 $T=691300 870360 1 0 $X=691300 $Y=864940
X2305 3970 3867 2 1 3990 3910 MUX2 $T=693160 769560 0 0 $X=693160 $Y=769180
X2306 3971 3956 2 1 4005 654 MUX2 $T=693160 830040 0 0 $X=693160 $Y=829660
X2307 3997 722 2 1 3968 681 MUX2 $T=698120 890520 1 180 $X=693780 $Y=890140
X2308 3980 3906 2 1 4010 3946 MUX2 $T=695020 749400 1 0 $X=695020 $Y=743980
X2309 4017 4009 2 1 4020 3609 MUX2 $T=700600 830040 0 0 $X=700600 $Y=829660
X2310 4049 4050 2 1 4021 3318 MUX2 $T=706180 870360 1 180 $X=701840 $Y=869980
X2311 4036 3822 2 1 4059 732 MUX2 $T=703700 739320 0 0 $X=703700 $Y=738940
X2312 4062 722 2 1 4025 728 MUX2 $T=708040 880440 0 180 $X=703700 $Y=875020
X2313 4038 685 2 1 734 732 MUX2 $T=704320 729240 1 0 $X=704320 $Y=723820
X2314 4043 3832 2 1 4064 4048 MUX2 $T=704940 809880 1 0 $X=704940 $Y=804460
X2315 3838 4050 2 1 4011 4057 MUX2 $T=711760 860280 0 180 $X=707420 $Y=854860
X2316 735 685 2 1 4087 3211 MUX2 $T=708040 739320 0 0 $X=708040 $Y=738940
X2317 4067 3867 2 1 4045 4048 MUX2 $T=708660 779640 1 0 $X=708660 $Y=774220
X2318 4094 3906 2 1 4073 732 MUX2 $T=713620 749400 1 180 $X=709280 $Y=749020
X2319 4074 3832 2 1 4116 3994 MUX2 $T=709280 809880 1 0 $X=709280 $Y=804460
X2320 4075 4009 2 1 4096 3994 MUX2 $T=709280 819960 1 0 $X=709280 $Y=814540
X2321 4083 3828 2 1 4108 4048 MUX2 $T=711140 789720 0 0 $X=711140 $Y=789340
X2322 4084 3828 2 1 4114 3994 MUX2 $T=711140 799800 0 0 $X=711140 $Y=799420
X2323 4026 754 2 1 4090 681 MUX2 $T=719200 890520 1 180 $X=714860 $Y=890140
X2324 758 757 2 1 750 3211 MUX2 $T=720440 729240 1 180 $X=716100 $Y=728860
X2325 4126 3947 2 1 4143 4130 MUX2 $T=717340 769560 0 0 $X=717340 $Y=769180
X2326 4145 3906 2 1 4128 4130 MUX2 $T=722300 749400 1 180 $X=717960 $Y=749020
X2327 4137 754 2 1 4154 752 MUX2 $T=719820 890520 0 0 $X=719820 $Y=890140
X2328 759 3867 2 1 4163 4130 MUX2 $T=721680 779640 1 0 $X=721680 $Y=774220
X2329 4157 4127 2 1 4168 4178 MUX2 $T=727260 819960 0 0 $X=727260 $Y=819580
X2330 4149 4159 2 1 4166 4198 MUX2 $T=729120 870360 1 0 $X=729120 $Y=864940
X2331 780 778 2 1 4216 752 MUX2 $T=732220 900600 1 0 $X=732220 $Y=895180
X2332 4259 804 2 1 4169 728 MUX2 $T=743380 890520 0 180 $X=739040 $Y=885100
X2333 800 4176 2 1 4171 4178 MUX2 $T=740900 819960 1 0 $X=740900 $Y=814540
X2334 801 778 2 1 4262 681 MUX2 $T=740900 900600 1 0 $X=740900 $Y=895180
X2335 4268 814 2 1 4194 4251 MUX2 $T=747100 749400 0 180 $X=742760 $Y=743980
X2336 4257 778 2 1 4277 728 MUX2 $T=744000 880440 0 0 $X=744000 $Y=880060
X2337 4260 4264 2 1 4291 4198 MUX2 $T=744620 870360 0 0 $X=744620 $Y=869980
X2338 4265 4234 2 1 4286 4178 MUX2 $T=745860 819960 1 0 $X=745860 $Y=814540
X2339 4270 4302 2 1 4274 768 MUX2 $T=753920 739320 1 180 $X=749580 $Y=738940
X2340 4306 4234 2 1 4342 4349 MUX2 $T=757640 840120 1 0 $X=757640 $Y=834700
X2341 4346 4352 2 1 4305 4178 MUX2 $T=763220 850200 1 180 $X=758880 $Y=849820
X2342 4377 4374 2 1 4301 4357 MUX2 $T=768180 850200 1 180 $X=763840 $Y=849820
X2343 4404 4360 2 1 4339 4381 MUX2 $T=772520 819960 0 180 $X=768180 $Y=814540
X2344 4406 4374 2 1 4351 4385 MUX2 $T=773140 850200 0 180 $X=768800 $Y=844780
X2345 4411 4407 2 1 4333 4381 MUX2 $T=773760 830040 1 180 $X=769420 $Y=829660
X2346 4349 4393 2 1 4320 873 MUX2 $T=782440 789720 1 180 $X=778100 $Y=789340
X2347 4451 4352 2 1 4465 4385 MUX2 $T=778100 850200 1 0 $X=778100 $Y=844780
X2348 4519 4505 2 1 4493 4349 MUX2 $T=790500 819960 0 180 $X=786160 $Y=814540
X2349 4508 4505 2 1 4494 4454 MUX2 $T=788640 809880 1 0 $X=788640 $Y=804460
X2350 4481 4512 2 1 4444 4454 MUX2 $T=789880 880440 0 0 $X=789880 $Y=880060
X2351 4523 4512 2 1 4542 4357 MUX2 $T=791120 850200 0 0 $X=791120 $Y=849820
X2352 4356 4560 2 1 4526 4349 MUX2 $T=796080 799800 0 180 $X=791740 $Y=794380
X2353 910 4560 2 1 4534 676 MUX2 $T=799180 830040 1 180 $X=794840 $Y=829660
X2354 4541 4505 2 1 4533 676 MUX2 $T=794840 840120 1 0 $X=794840 $Y=834700
X2355 4632 4539 2 1 4559 888 MUX2 $T=806000 779640 1 180 $X=801660 $Y=779260
X2356 4622 4585 2 1 4586 923 MUX2 $T=810960 749400 1 180 $X=806620 $Y=749020
X2357 4651 4505 2 1 4673 4381 MUX2 $T=811580 809880 0 0 $X=811580 $Y=809500
X2358 4669 4539 2 1 4690 4687 MUX2 $T=814680 779640 0 0 $X=814680 $Y=779260
X2359 4594 4407 2 1 4693 4717 MUX2 $T=815300 819960 1 0 $X=815300 $Y=814540
X2360 4722 4608 2 1 4679 4687 MUX2 $T=823360 779640 1 180 $X=819020 $Y=779260
X2361 4599 4702 2 1 4715 4676 MUX2 $T=819020 850200 1 0 $X=819020 $Y=844780
X2362 4747 4699 2 1 4682 923 MUX2 $T=825220 749400 0 180 $X=820880 $Y=743980
X2363 4694 4731 2 1 4640 4676 MUX2 $T=827080 830040 1 180 $X=822740 $Y=829660
X2364 4759 4585 2 1 4678 4740 MUX2 $T=830800 759480 0 180 $X=826460 $Y=754060
X2365 4762 4702 2 1 4742 4717 MUX2 $T=830800 840120 0 180 $X=826460 $Y=834700
X2366 4654 4608 2 1 4745 4740 MUX2 $T=831420 789720 0 180 $X=827080 $Y=784300
X2367 4548 4731 2 1 4729 4717 MUX2 $T=831420 830040 1 180 $X=827080 $Y=829660
X2368 4750 4699 2 1 4767 4740 MUX2 $T=828320 749400 1 0 $X=828320 $Y=743980
X2369 4770 4575 2 1 4733 4740 MUX2 $T=832660 769560 0 180 $X=828320 $Y=764140
X2370 4776 4645 2 1 4709 952 MUX2 $T=833280 729240 0 180 $X=828940 $Y=723820
X2371 4724 4785 2 1 4765 4740 MUX2 $T=835140 799800 1 180 $X=830800 $Y=799420
X2372 4331 4645 2 1 956 959 MUX2 $T=831420 729240 0 0 $X=831420 $Y=728860
X2373 4579 4450 2 1 4718 4717 MUX2 $T=838240 819960 0 180 $X=833900 $Y=814540
X2374 4794 4814 2 1 4696 4717 MUX2 $T=838860 830040 1 180 $X=834520 $Y=829660
X2375 4803 4822 2 1 4793 4717 MUX2 $T=839480 830040 0 180 $X=835140 $Y=824620
X2376 4827 4699 2 1 4799 4687 MUX2 $T=841340 739320 1 180 $X=837000 $Y=738940
X2377 4841 4575 2 1 4809 4819 MUX2 $T=845060 759480 1 180 $X=840720 $Y=759100
X2378 4816 4820 2 1 4844 4819 MUX2 $T=840720 779640 0 0 $X=840720 $Y=779260
X2379 4845 4785 2 1 4811 4819 MUX2 $T=846300 799800 1 180 $X=841960 $Y=799420
X2380 4828 4450 2 1 4851 4819 MUX2 $T=841960 819960 1 0 $X=841960 $Y=814540
X2381 4843 4822 2 1 4823 4676 MUX2 $T=846300 840120 0 180 $X=841960 $Y=834700
X2382 4829 4585 2 1 4861 4819 MUX2 $T=842580 759480 1 0 $X=842580 $Y=754060
X2383 4853 4801 2 1 4796 4819 MUX2 $T=846920 789720 0 180 $X=842580 $Y=784300
X2384 4834 960 2 1 4862 4687 MUX2 $T=843820 739320 1 0 $X=843820 $Y=733900
X2385 4644 4814 2 1 4868 4676 MUX2 $T=846300 840120 1 0 $X=846300 $Y=834700
X2386 4881 4837 2 1 4864 4676 MUX2 $T=853740 819960 1 180 $X=849400 $Y=819580
X2387 4909 4777 2 1 4865 4888 MUX2 $T=857460 789720 0 180 $X=853120 $Y=784300
X2388 4923 4887 2 1 4885 4687 MUX2 $T=860560 739320 1 180 $X=856220 $Y=738940
X2389 4924 4903 2 1 4905 4687 MUX2 $T=860560 759480 0 180 $X=856220 $Y=754060
X2390 983 4903 2 1 4894 4888 MUX2 $T=862420 769560 0 180 $X=858080 $Y=764140
X2391 4935 4801 2 1 4886 4888 MUX2 $T=862420 789720 0 180 $X=858080 $Y=784300
X2392 4925 4785 2 1 4896 3910 MUX2 $T=863040 799800 1 180 $X=858700 $Y=799420
X2393 4939 4910 2 1 4921 4385 MUX2 $T=864280 860280 0 180 $X=859940 $Y=854860
X2394 4920 4887 2 1 4940 4899 MUX2 $T=860560 739320 0 0 $X=860560 $Y=738940
X2395 4946 4882 2 1 4917 4901 MUX2 $T=864900 890520 0 180 $X=860560 $Y=885100
X2396 4664 4785 2 1 4855 4953 MUX2 $T=862420 799800 1 0 $X=862420 $Y=794380
X2397 4787 4830 2 1 4954 4385 MUX2 $T=862420 840120 1 0 $X=862420 $Y=834700
X2398 4941 4897 2 1 4944 4385 MUX2 $T=869240 850200 1 180 $X=864900 $Y=849820
X2399 4904 4785 2 1 4880 4975 MUX2 $T=866140 809880 0 0 $X=866140 $Y=809500
X2400 4990 4887 2 1 4967 924 MUX2 $T=873580 749400 1 180 $X=869240 $Y=749020
X2401 4949 4777 2 1 5001 5008 MUX2 $T=869240 779640 1 0 $X=869240 $Y=774220
X2402 4958 4801 2 1 4928 4953 MUX2 $T=874820 789720 1 180 $X=870480 $Y=789340
X2403 4998 4801 2 1 4966 4975 MUX2 $T=874820 809880 1 180 $X=870480 $Y=809500
X2404 5013 960 2 1 4987 639 MUX2 $T=876680 739320 0 180 $X=872340 $Y=733900
X2405 5002 4903 2 1 4971 4953 MUX2 $T=876680 759480 1 180 $X=872340 $Y=759100
X2406 4999 985 2 1 4986 991 MUX2 $T=876680 890520 0 180 $X=872340 $Y=885100
X2407 4984 985 2 1 994 992 MUX2 $T=876680 890520 1 180 $X=872340 $Y=890140
X2408 4996 4830 2 1 4989 5016 MUX2 $T=873580 840120 1 0 $X=873580 $Y=834700
X2409 999 964 2 1 995 639 MUX2 $T=878540 729240 0 180 $X=874200 $Y=723820
X2410 5027 4820 2 1 5063 4888 MUX2 $T=879780 779640 1 0 $X=879780 $Y=774220
X2411 5028 4916 2 1 5051 4970 MUX2 $T=879780 870360 0 0 $X=879780 $Y=869980
X2412 5066 4820 2 1 5014 5008 MUX2 $T=885360 789720 1 180 $X=881020 $Y=789340
X2413 5040 4837 2 1 4978 4888 MUX2 $T=882260 819960 1 0 $X=882260 $Y=814540
X2414 5071 4887 2 1 5045 5010 MUX2 $T=887220 759480 1 180 $X=882880 $Y=759100
X2415 4983 4887 2 1 5007 1014 MUX2 $T=883500 739320 1 0 $X=883500 $Y=733900
X2416 5035 4821 2 1 5054 4953 MUX2 $T=889080 799800 0 180 $X=884740 $Y=794380
X2417 5029 938 2 1 5085 992 MUX2 $T=884740 900600 1 0 $X=884740 $Y=895180
X2418 5092 4821 2 1 5050 4975 MUX2 $T=890940 819960 0 180 $X=886600 $Y=814540
X2419 5072 4830 2 1 5094 5096 MUX2 $T=886600 840120 0 0 $X=886600 $Y=839740
X2420 5074 4830 2 1 4985 5095 MUX2 $T=886600 860280 0 0 $X=886600 $Y=859900
X2421 5079 4887 2 1 5097 1018 MUX2 $T=887840 739320 1 0 $X=887840 $Y=733900
X2422 1023 4821 2 1 5099 4888 MUX2 $T=895900 799800 0 180 $X=891560 $Y=794380
X2423 5125 4821 2 1 5104 5010 MUX2 $T=896520 809880 1 180 $X=892180 $Y=809500
X2424 5105 4916 2 1 5126 5095 MUX2 $T=892180 860280 0 0 $X=892180 $Y=859900
X2425 5075 938 2 1 5133 991 MUX2 $T=892180 890520 0 0 $X=892180 $Y=890140
X2426 5068 4897 2 1 5076 5016 MUX2 $T=899000 840120 0 180 $X=894660 $Y=834700
X2427 5118 4916 2 1 5135 1020 MUX2 $T=894660 870360 0 0 $X=894660 $Y=869980
X2428 1028 960 2 1 5123 1025 MUX2 $T=900240 729240 0 180 $X=895900 $Y=723820
X2429 5124 4820 2 1 5143 1026 MUX2 $T=895900 789720 0 0 $X=895900 $Y=789340
X2430 5127 4903 2 1 5158 1018 MUX2 $T=897140 749400 0 0 $X=897140 $Y=749020
X2431 1027 4903 2 1 5161 5010 MUX2 $T=897760 759480 0 0 $X=897760 $Y=759100
X2432 5139 4897 2 1 5167 5096 MUX2 $T=899620 840120 1 0 $X=899620 $Y=834700
X2433 5148 964 2 1 5171 1018 MUX2 $T=900860 729240 1 0 $X=900860 $Y=723820
X2434 5156 4897 2 1 5182 5095 MUX2 $T=901480 850200 0 0 $X=901480 $Y=849820
X2435 5163 4820 2 1 5082 5179 MUX2 $T=902720 779640 1 0 $X=902720 $Y=774220
X2436 5164 4821 2 1 5198 1018 MUX2 $T=902720 799800 1 0 $X=902720 $Y=794380
X2437 5187 4910 2 1 5110 4970 MUX2 $T=907060 870360 1 180 $X=902720 $Y=869980
X2438 1033 1030 2 1 5196 991 MUX2 $T=904580 890520 0 0 $X=904580 $Y=890140
X2439 5146 960 2 1 5201 5179 MUX2 $T=905820 739320 1 0 $X=905820 $Y=733900
X2440 5205 4837 2 1 5184 5183 MUX2 $T=910780 819960 0 180 $X=906440 $Y=814540
X2441 5186 4910 2 1 5213 5016 MUX2 $T=906440 840120 0 0 $X=906440 $Y=839740
X2442 5188 4910 2 1 5206 1020 MUX2 $T=906440 880440 0 0 $X=906440 $Y=880060
X2443 5190 4897 2 1 5207 4970 MUX2 $T=907060 870360 0 0 $X=907060 $Y=869980
X2444 5204 4837 2 1 5215 1026 MUX2 $T=910160 809880 0 0 $X=910160 $Y=809500
X2445 5208 4820 2 1 5222 5195 MUX2 $T=911400 789720 1 0 $X=911400 $Y=784300
X2446 5209 4837 2 1 5229 5185 MUX2 $T=911400 809880 1 0 $X=911400 $Y=804460
X2447 5210 4897 2 1 5218 1020 MUX2 $T=911400 870360 0 0 $X=911400 $Y=869980
X2448 5220 4837 2 1 5239 5195 MUX2 $T=915120 809880 0 0 $X=915120 $Y=809500
X2449 5243 5233 2 1 5200 5221 MUX2 $T=920080 769560 1 180 $X=915740 $Y=769180
X2450 5259 5212 2 1 5197 1046 MUX2 $T=924420 749400 1 180 $X=920080 $Y=749020
X2451 5273 5286 2 1 5249 1046 MUX2 $T=928140 739320 0 180 $X=923800 $Y=733900
X2452 5276 5267 2 1 5238 5221 MUX2 $T=928140 779640 0 180 $X=923800 $Y=774220
X2453 5277 5269 2 1 5223 5261 MUX2 $T=928140 870360 0 180 $X=923800 $Y=864940
X2454 5279 5280 2 1 5228 1046 MUX2 $T=928760 749400 1 180 $X=924420 $Y=749020
X2455 5282 5260 2 1 5236 5221 MUX2 $T=928760 799800 0 180 $X=924420 $Y=794380
X2456 5290 5285 2 1 5230 5185 MUX2 $T=930000 819960 1 180 $X=925660 $Y=819580
X2457 5232 5291 2 1 5254 991 MUX2 $T=930000 850200 0 180 $X=925660 $Y=844780
X2458 1052 5269 2 1 5224 1048 MUX2 $T=931860 870360 1 180 $X=927520 $Y=869980
X2459 5313 5297 2 1 5251 1048 MUX2 $T=931860 880440 1 180 $X=927520 $Y=880060
X2460 5281 5267 2 1 5314 5261 MUX2 $T=928140 779640 1 0 $X=928140 $Y=774220
X2461 5322 5323 2 1 5258 5185 MUX2 $T=934340 819960 1 180 $X=930000 $Y=819580
X2462 5339 5280 2 1 5246 5179 MUX2 $T=937440 759480 1 180 $X=933100 $Y=759100
X2463 5341 5338 2 1 5271 5179 MUX2 $T=938060 749400 1 180 $X=933720 $Y=749020
X2464 5349 5291 2 1 5292 4976 MUX2 $T=938060 850200 0 180 $X=933720 $Y=844780
X2465 5351 1057 2 1 5240 1053 MUX2 $T=938680 900600 0 180 $X=934340 $Y=895180
X2466 5352 5345 2 1 5306 5221 MUX2 $T=939300 789720 1 180 $X=934960 $Y=789340
X2467 5353 5260 2 1 5315 5261 MUX2 $T=939300 799800 0 180 $X=934960 $Y=794380
X2468 5357 5286 2 1 5300 1054 MUX2 $T=939920 739320 1 180 $X=935580 $Y=738940
X2469 5365 5330 2 1 5327 5261 MUX2 $T=941160 779640 1 180 $X=936820 $Y=779260
X2470 5376 1055 2 1 1059 1054 MUX2 $T=942400 729240 0 180 $X=938060 $Y=723820
X2471 5344 5280 2 1 5368 1064 MUX2 $T=938060 749400 0 0 $X=938060 $Y=749020
X2472 5346 5345 2 1 5343 5261 MUX2 $T=943020 809880 0 180 $X=938680 $Y=804460
X2473 5390 5304 2 1 5336 5234 MUX2 $T=944260 880440 0 180 $X=939920 $Y=875020
X2474 5388 5256 2 1 5334 5354 MUX2 $T=946120 840120 1 180 $X=941780 $Y=839740
X2475 5399 5291 2 1 5272 5354 MUX2 $T=947360 860280 1 180 $X=943020 $Y=859900
X2476 5383 5345 2 1 5408 5354 MUX2 $T=943640 809880 1 0 $X=943640 $Y=804460
X2477 5387 5330 2 1 5414 5354 MUX2 $T=944260 789720 0 0 $X=944260 $Y=789340
X2478 5398 5323 2 1 5433 5354 MUX2 $T=946740 850200 0 0 $X=946740 $Y=849820
X2479 1073 5434 2 1 5402 5234 MUX2 $T=951080 890520 1 180 $X=946740 $Y=890140
X2480 5409 5285 2 1 5429 1074 MUX2 $T=947360 819960 0 0 $X=947360 $Y=819580
X2481 5419 1055 2 1 1077 1035 MUX2 $T=948600 729240 1 0 $X=948600 $Y=723820
X2482 5441 5325 2 1 5423 5234 MUX2 $T=953560 880440 0 180 $X=949220 $Y=875020
X2483 5455 5285 2 1 5430 5354 MUX2 $T=955420 870360 1 180 $X=951080 $Y=869980
X2484 5463 5323 2 1 5389 1074 MUX2 $T=956660 819960 0 180 $X=952320 $Y=814540
X2485 5436 5434 2 1 5464 5195 MUX2 $T=952320 840120 0 0 $X=952320 $Y=839740
X2486 5476 1075 2 1 5443 4901 MUX2 $T=957900 890520 0 180 $X=953560 $Y=885100
X2487 5470 5323 2 1 5489 5195 MUX2 $T=956660 819960 1 0 $X=956660 $Y=814540
X2488 5490 5291 2 1 5467 5195 MUX2 $T=961000 840120 1 180 $X=956660 $Y=839740
X2489 5493 5393 2 1 5506 1071 MUX2 $T=961000 739320 1 0 $X=961000 $Y=733900
X2490 1088 1057 2 1 5487 5497 MUX2 $T=965340 890520 0 180 $X=961000 $Y=885100
X2491 5498 1055 2 1 1089 1071 MUX2 $T=961620 729240 1 0 $X=961620 $Y=723820
X2492 5502 5338 2 1 5520 1071 MUX2 $T=962860 759480 1 0 $X=962860 $Y=754060
X2493 5491 5434 2 1 5505 5183 MUX2 $T=967820 840120 1 180 $X=963480 $Y=839740
X2494 1091 1055 2 1 1094 1080 MUX2 $T=966580 729240 1 0 $X=966580 $Y=723820
X2495 5521 5330 2 1 5566 5557 MUX2 $T=966580 789720 1 0 $X=966580 $Y=784300
X2496 5556 5304 2 1 5533 5497 MUX2 $T=972160 860280 1 180 $X=967820 $Y=859900
X2497 5544 5345 2 1 5593 5557 MUX2 $T=970300 789720 0 0 $X=970300 $Y=789340
X2498 5545 5323 2 1 5570 5183 MUX2 $T=970300 819960 0 0 $X=970300 $Y=819580
X2499 5546 5291 2 1 5571 5183 MUX2 $T=970300 850200 1 0 $X=970300 $Y=844780
X2500 5549 1055 2 1 5574 1098 MUX2 $T=970920 729240 1 0 $X=970920 $Y=723820
X2501 5486 5403 2 1 5529 5497 MUX2 $T=976500 759480 1 180 $X=972160 $Y=759100
X2502 5586 1075 2 1 5531 5497 MUX2 $T=976500 890520 0 180 $X=972160 $Y=885100
X2503 5576 5427 2 1 5619 1097 MUX2 $T=975260 779640 1 0 $X=975260 $Y=774220
X2504 5613 5325 2 1 5592 5557 MUX2 $T=980840 880440 0 180 $X=976500 $Y=875020
X2505 5595 5403 2 1 5615 1074 MUX2 $T=977120 769560 1 0 $X=977120 $Y=764140
X2506 5597 5291 2 1 5634 5600 MUX2 $T=977120 850200 1 0 $X=977120 $Y=844780
X2507 1101 1075 2 1 1106 1105 MUX2 $T=977120 900600 1 0 $X=977120 $Y=895180
X2508 5604 5338 2 1 5624 1074 MUX2 $T=978980 749400 1 0 $X=978980 $Y=743980
X2509 5609 5323 2 1 5630 5600 MUX2 $T=979600 830040 1 0 $X=979600 $Y=824620
X2510 5610 5285 2 1 5632 5600 MUX2 $T=979600 840120 1 0 $X=979600 $Y=834700
X2511 5617 5434 2 1 5642 5600 MUX2 $T=980840 840120 0 0 $X=980840 $Y=839740
X2512 5618 5325 2 1 5633 5497 MUX2 $T=980840 880440 1 0 $X=980840 $Y=875020
X2513 5620 5393 2 1 5636 1098 MUX2 $T=981460 739320 1 0 $X=981460 $Y=733900
X2514 5626 5403 2 1 5646 5600 MUX2 $T=982700 759480 0 0 $X=982700 $Y=759100
X2515 5684 5666 2 1 5623 1105 MUX2 $T=998820 890520 1 180 $X=994480 $Y=890140
X2516 5728 5724 2 1 5629 1105 MUX2 $T=1003160 890520 1 180 $X=998820 $Y=890140
X2517 5740 5733 2 1 5643 1097 MUX2 $T=1005020 789720 0 180 $X=1000680 $Y=784300
X2518 5759 5720 2 1 5725 1097 MUX2 $T=1007500 769560 0 180 $X=1003160 $Y=764140
X2519 5776 5700 2 1 5712 1097 MUX2 $T=1011220 759480 1 180 $X=1006880 $Y=759100
X2520 5898 5802 2 1 5977 5956 MUX2 $T=1050900 830040 1 180 $X=1046560 $Y=829660
X2521 5971 5794 2 1 6005 1185 MUX2 $T=1046560 880440 1 0 $X=1046560 $Y=875020
X2522 5999 5863 2 1 6019 6018 MUX2 $T=1050280 759480 1 0 $X=1050280 $Y=754060
X2523 6025 5666 2 1 5978 1185 MUX2 $T=1054620 880440 1 180 $X=1050280 $Y=880060
X2524 6014 5955 2 1 6021 6018 MUX2 $T=1059580 809880 1 180 $X=1055240 $Y=809500
X2525 6030 6024 2 1 6038 6047 MUX2 $T=1055240 860280 1 0 $X=1055240 $Y=854860
X2526 6051 5888 2 1 6009 6018 MUX2 $T=1061440 779640 1 180 $X=1057100 $Y=779260
X2527 6057 5910 2 1 6035 6018 MUX2 $T=1061440 789720 1 180 $X=1057100 $Y=789340
X2528 6042 6041 2 1 6059 6047 MUX2 $T=1058340 870360 0 0 $X=1058340 $Y=869980
X2529 6070 6048 2 1 6043 6047 MUX2 $T=1063300 850200 0 180 $X=1058960 $Y=844780
X2530 6052 5900 2 1 6066 6018 MUX2 $T=1059580 809880 0 0 $X=1059580 $Y=809500
X2531 6040 1195 2 1 6007 6047 MUX2 $T=1064540 890520 1 180 $X=1060200 $Y=890140
X2532 6061 6026 2 1 6034 6065 MUX2 $T=1067020 830040 0 180 $X=1062680 $Y=824620
X2533 6086 6036 2 1 6044 6047 MUX2 $T=1067020 870360 1 180 $X=1062680 $Y=869980
X2534 6105 6020 2 1 6029 6065 MUX2 $T=1070740 819960 1 180 $X=1066400 $Y=819580
X2535 6089 6093 2 1 6112 6098 MUX2 $T=1067640 779640 1 0 $X=1067640 $Y=774220
X2536 1203 1202 2 1 6074 1199 MUX2 $T=1072600 729240 1 180 $X=1068260 $Y=728860
X2537 6118 6091 2 1 6097 6098 MUX2 $T=1073840 749400 1 180 $X=1069500 $Y=749020
X2538 6119 6048 2 1 6101 6102 MUX2 $T=1073840 850200 1 180 $X=1069500 $Y=849820
X2539 6126 6104 2 1 6087 6107 MUX2 $T=1075080 809880 0 180 $X=1070740 $Y=804460
X2540 6076 6084 2 1 6132 6098 MUX2 $T=1071980 779640 1 0 $X=1071980 $Y=774220
X2541 6113 6020 2 1 6115 6107 MUX2 $T=1076320 830040 0 180 $X=1071980 $Y=824620
X2542 1204 1194 2 1 1210 6122 MUX2 $T=1072600 729240 1 0 $X=1072600 $Y=723820
X2543 6121 6091 2 1 6137 6122 MUX2 $T=1073840 759480 1 0 $X=1073840 $Y=754060
X2544 6143 6104 2 1 6117 5581 MUX2 $T=1079420 809880 1 180 $X=1075080 $Y=809500
X2545 6144 6036 2 1 6083 6102 MUX2 $T=1079420 870360 0 180 $X=1075080 $Y=864940
X2546 1215 6024 2 1 6111 6102 MUX2 $T=1079420 880440 0 180 $X=1075080 $Y=875020
X2547 1206 1208 2 1 1218 6148 MUX2 $T=1075700 900600 1 0 $X=1075700 $Y=895180
X2548 6134 6093 2 1 6141 6122 MUX2 $T=1076320 779640 1 0 $X=1076320 $Y=774220
X2549 6155 6026 2 1 6131 6107 MUX2 $T=1080660 830040 0 180 $X=1076320 $Y=824620
X2550 1211 1202 2 1 6152 6122 MUX2 $T=1076940 729240 1 0 $X=1076940 $Y=723820
X2551 6170 6084 2 1 6130 6122 MUX2 $T=1083760 779640 1 180 $X=1079420 $Y=779260
X2552 1217 1205 2 1 6167 6102 MUX2 $T=1079420 890520 0 0 $X=1079420 $Y=890140
X2553 6142 6153 2 1 6114 6122 MUX2 $T=1085000 759480 0 180 $X=1080660 $Y=754060
X2554 6154 6082 2 1 6181 5581 MUX2 $T=1080660 799800 0 0 $X=1080660 $Y=799420
X2555 6177 1194 2 1 1219 1220 MUX2 $T=1085620 729240 0 180 $X=1081280 $Y=723820
X2556 6192 6048 2 1 6158 6148 MUX2 $T=1088100 850200 1 180 $X=1083760 $Y=849820
X2557 6173 6041 2 1 6198 6102 MUX2 $T=1084380 870360 1 0 $X=1084380 $Y=864940
X2558 6203 6082 2 1 6182 6098 MUX2 $T=1090580 809880 0 180 $X=1086240 $Y=804460
X2559 6175 6093 2 1 6219 6107 MUX2 $T=1087480 789720 0 0 $X=1087480 $Y=789340
X2560 6191 6091 2 1 6214 1220 MUX2 $T=1089340 749400 0 0 $X=1089340 $Y=749020
X2561 6233 6020 2 1 6200 5581 MUX2 $T=1095540 830040 0 180 $X=1091200 $Y=824620
X2562 6236 6084 2 1 6212 1220 MUX2 $T=1096780 779640 0 180 $X=1092440 $Y=774220
X2563 6240 6082 2 1 6208 6107 MUX2 $T=1097400 809880 0 180 $X=1093060 $Y=804460
X2564 6222 6036 2 1 6245 1230 MUX2 $T=1093060 880440 1 0 $X=1093060 $Y=875020
X2565 1233 1202 2 1 6213 1220 MUX2 $T=1098640 729240 0 180 $X=1094300 $Y=723820
X2566 6252 6026 2 1 6215 6226 MUX2 $T=1098640 840120 0 180 $X=1094300 $Y=834700
X2567 6229 6036 2 1 6257 6148 MUX2 $T=1094920 880440 0 0 $X=1094920 $Y=880060
X2568 6247 6041 2 1 6268 1230 MUX2 $T=1098020 880440 1 0 $X=1098020 $Y=875020
X2569 6258 6082 2 1 6274 6273 MUX2 $T=1099880 809880 1 0 $X=1099880 $Y=804460
X2570 6265 6153 2 1 6283 1238 MUX2 $T=1101740 749400 0 0 $X=1101740 $Y=749020
X2571 6266 6020 2 1 6288 6226 MUX2 $T=1101740 830040 1 0 $X=1101740 $Y=824620
X2572 6289 6048 2 1 6264 1230 MUX2 $T=1106080 850200 1 180 $X=1101740 $Y=849820
X2573 6292 1202 2 1 6230 1209 MUX2 $T=1106700 729240 0 180 $X=1102360 $Y=723820
X2574 6272 6084 2 1 6291 6293 MUX2 $T=1102980 779640 1 0 $X=1102980 $Y=774220
X2575 6277 6093 2 1 6314 6273 MUX2 $T=1104220 789720 0 0 $X=1104220 $Y=789340
X2576 6295 6020 2 1 6318 6273 MUX2 $T=1106080 830040 1 0 $X=1106080 $Y=824620
X2577 6300 6024 2 1 6321 1230 MUX2 $T=1106700 850200 0 0 $X=1106700 $Y=849820
X2578 6301 6091 2 1 6279 1238 MUX2 $T=1107320 739320 0 0 $X=1107320 $Y=738940
X2579 6309 6104 2 1 6346 6065 MUX2 $T=1108560 809880 0 0 $X=1108560 $Y=809500
X2580 6344 6036 2 1 6276 1243 MUX2 $T=1112900 890520 1 180 $X=1108560 $Y=890140
X2581 6320 6020 2 1 6349 6081 MUX2 $T=1110420 830040 1 0 $X=1110420 $Y=824620
X2582 6330 6048 2 1 6350 1251 MUX2 $T=1111660 850200 0 0 $X=1111660 $Y=849820
X2583 6353 1202 2 1 6332 1238 MUX2 $T=1116620 739320 0 180 $X=1112280 $Y=733900
X2584 6333 6091 2 1 6354 1252 MUX2 $T=1112280 739320 0 0 $X=1112280 $Y=738940
X2585 6334 6153 2 1 6355 1252 MUX2 $T=1112280 749400 0 0 $X=1112280 $Y=749020
X2586 6335 6153 2 1 6356 6293 MUX2 $T=1112280 759480 1 0 $X=1112280 $Y=754060
X2587 6336 6084 2 1 6357 1238 MUX2 $T=1112280 759480 0 0 $X=1112280 $Y=759100
X2588 6244 6093 2 1 6358 1187 MUX2 $T=1112280 779640 0 0 $X=1112280 $Y=779260
X2589 6331 6026 2 1 6359 6081 MUX2 $T=1112280 840120 1 0 $X=1112280 $Y=834700
X2590 1249 6024 2 1 6360 1251 MUX2 $T=1112280 860280 0 0 $X=1112280 $Y=859900
X2591 6342 6082 2 1 6365 1187 MUX2 $T=1112900 799800 0 0 $X=1112900 $Y=799420
X2592 6343 6082 2 1 6366 6065 MUX2 $T=1112900 809880 1 0 $X=1112900 $Y=804460
X2593 6345 1202 2 1 6368 1252 MUX2 $T=1114140 729240 1 0 $X=1114140 $Y=723820
X2594 6351 6041 2 1 6363 1251 MUX2 $T=1120340 880440 1 180 $X=1116000 $Y=880060
X2595 6370 6048 2 1 6373 6081 MUX2 $T=1120340 850200 1 0 $X=1120340 $Y=844780
X2596 6371 6041 2 1 6372 6081 MUX2 $T=1120340 880440 0 0 $X=1120340 $Y=880060
X2597 1370 14 1375 1398 1 18 2 AOI22S $T=230640 729240 1 0 $X=230640 $Y=723820
X2598 1370 26 1465 28 1 31 2 AOI22S $T=243660 729240 1 0 $X=243660 $Y=723820
X2599 1453 1599 1594 37 1 1580 2 AOI22S $T=264740 860280 0 0 $X=264740 $Y=859900
X2600 1856 127 1659 1855 1 144 2 AOI22S $T=313100 860280 0 0 $X=313100 $Y=859900
X2601 145 139 1821 149 1 132 2 AOI22S $T=316200 890520 1 0 $X=316200 $Y=885100
X2602 74 168 1951 161 1 132 2 AOI22S $T=330460 900600 0 180 $X=326740 $Y=895180
X2603 2156 2177 2142 2161 1 217 2 AOI22S $T=362080 870360 0 0 $X=362080 $Y=869980
X2604 2311 2330 2412 2211 1 2420 2 AOI22S $T=398660 870360 0 0 $X=398660 $Y=869980
X2605 2689 2674 2683 2639 1 2559 2 AOI22S $T=448880 799800 0 180 $X=445160 $Y=794380
X2606 2689 2674 2677 2619 1 2597 2 AOI22S $T=450120 789720 1 180 $X=446400 $Y=789340
X2607 2700 2690 2693 2602 1 2427 2 AOI22S $T=450120 830040 1 180 $X=446400 $Y=829660
X2608 359 355 2732 2676 1 2552 2 AOI22S $T=457560 890520 0 180 $X=453840 $Y=885100
X2609 2689 2674 2733 2598 1 2724 2 AOI22S $T=458180 799800 0 180 $X=454460 $Y=794380
X2610 2700 2690 2743 2709 1 2499 2 AOI22S $T=460660 830040 1 180 $X=456940 $Y=829660
X2611 359 355 2750 2741 1 2740 2 AOI22S $T=461900 890520 0 180 $X=458180 $Y=885100
X2612 2756 361 2754 2746 1 2721 2 AOI22S $T=462520 880440 0 180 $X=458800 $Y=875020
X2613 2700 2690 2765 2628 1 2565 2 AOI22S $T=464380 830040 1 180 $X=460660 $Y=829660
X2614 2689 2739 2783 2759 1 2744 2 AOI22S $T=467480 799800 0 180 $X=463760 $Y=794380
X2615 2689 2739 2780 2543 1 2627 2 AOI22S $T=465620 789720 0 0 $X=465620 $Y=789340
X2616 2700 2690 2805 2827 1 2804 2 AOI22S $T=471820 840120 1 0 $X=471820 $Y=834700
X2617 2689 2739 2858 2811 1 2668 2 AOI22S $T=479260 799800 0 180 $X=475540 $Y=794380
X2618 2700 2843 2855 2850 1 2835 2 AOI22S $T=481740 830040 1 180 $X=478020 $Y=829660
X2619 396 391 2853 2757 1 390 2 AOI22S $T=485460 900600 0 180 $X=481740 $Y=895180
X2620 2895 391 2885 2355 1 388 2 AOI22S $T=488560 870360 0 180 $X=484840 $Y=864940
X2621 2895 361 2894 2880 1 2859 2 AOI22S $T=489180 860280 1 180 $X=485460 $Y=859900
X2622 2756 2843 2903 2840 1 2889 2 AOI22S $T=491040 830040 0 180 $X=487320 $Y=824620
X2623 396 391 2896 2886 1 2908 2 AOI22S $T=487940 880440 0 0 $X=487940 $Y=880060
X2624 2879 2739 2915 2924 1 2411 2 AOI22S $T=492280 799800 0 0 $X=492280 $Y=799420
X2625 2951 2931 2936 2861 1 400 2 AOI22S $T=499100 749400 1 180 $X=495380 $Y=749020
X2626 2756 2843 2919 2899 1 2943 2 AOI22S $T=496000 830040 0 0 $X=496000 $Y=829660
X2627 2951 2931 2957 2822 1 2934 2 AOI22S $T=500340 759480 0 180 $X=496620 $Y=754060
X2628 2951 2931 2960 2916 1 407 2 AOI22S $T=502820 749400 1 180 $X=499100 $Y=749020
X2629 2951 2931 2970 2792 1 406 2 AOI22S $T=504680 749400 0 180 $X=500960 $Y=743980
X2630 423 2929 2980 412 1 410 2 AOI22S $T=504680 900600 0 180 $X=500960 $Y=895180
X2631 2756 2843 2974 2920 1 2992 2 AOI22S $T=503440 830040 0 0 $X=503440 $Y=829660
X2632 396 391 2990 2550 1 3001 2 AOI22S $T=505300 880440 0 0 $X=505300 $Y=880060
X2633 2951 2931 3026 3009 1 2981 2 AOI22S $T=511500 769560 0 180 $X=507780 $Y=764140
X2634 423 2929 3008 3013 1 408 2 AOI22S $T=508400 900600 1 0 $X=508400 $Y=895180
X2635 2879 3054 3057 3027 1 3048 2 AOI22S $T=520800 799800 1 180 $X=517080 $Y=799420
X2636 3077 355 3067 2251 1 3051 2 AOI22S $T=522660 870360 0 180 $X=518940 $Y=864940
X2637 3053 3021 3066 3037 1 3029 2 AOI22S $T=523900 819960 1 180 $X=520180 $Y=819580
X2638 3099 3084 3069 3071 1 3059 2 AOI22S $T=528240 759480 1 180 $X=524520 $Y=759100
X2639 3077 3054 3100 3114 1 3088 2 AOI22S $T=526380 799800 1 0 $X=526380 $Y=794380
X2640 3053 3021 3113 3122 1 3105 2 AOI22S $T=527620 819960 0 0 $X=527620 $Y=819580
X2641 423 420 3111 441 1 442 2 AOI22S $T=528240 900600 1 0 $X=528240 $Y=895180
X2642 3077 3054 3124 2383 1 2989 2 AOI22S $T=528860 809880 1 0 $X=528860 $Y=804460
X2643 3053 3021 3127 3132 1 2398 2 AOI22S $T=530100 860280 1 0 $X=530100 $Y=854860
X2644 3053 3021 3115 3139 1 3126 2 AOI22S $T=530720 850200 0 0 $X=530720 $Y=849820
X2645 3053 429 3136 3129 1 3147 2 AOI22S $T=531340 819960 0 0 $X=531340 $Y=819580
X2646 3099 3084 3043 3160 1 3154 2 AOI22S $T=533820 759480 0 0 $X=533820 $Y=759100
X2647 3099 3084 3207 462 1 3170 2 AOI22S $T=545600 759480 0 0 $X=545600 $Y=759100
X2648 3035 3045 3228 3219 1 3182 2 AOI22S $T=550560 769560 0 0 $X=550560 $Y=769180
X2649 3280 3262 3274 3235 1 3222 2 AOI22S $T=561100 819960 0 180 $X=557380 $Y=814540
X2650 3210 3202 3254 3273 1 3279 2 AOI22S $T=558000 749400 0 0 $X=558000 $Y=749020
X2651 3280 3262 3281 3266 1 3184 2 AOI22S $T=561720 840120 1 180 $X=558000 $Y=839740
X2652 3035 3045 3272 3206 1 3292 2 AOI22S $T=559240 779640 1 0 $X=559240 $Y=774220
X2653 3298 3045 3300 3276 1 3176 2 AOI22S $T=563580 769560 1 180 $X=559860 $Y=769180
X2654 486 3297 3302 3242 1 3218 2 AOI22S $T=565440 880440 1 180 $X=561720 $Y=880060
X2655 3330 3297 3348 3289 1 3278 2 AOI22S $T=569780 850200 0 180 $X=566060 $Y=844780
X2656 3330 3297 3329 3214 1 3249 2 AOI22S $T=571020 860280 0 180 $X=567300 $Y=854860
X2657 486 493 3341 492 1 479 2 AOI22S $T=571020 900600 0 180 $X=567300 $Y=895180
X2658 486 3297 3331 2493 1 470 2 AOI22S $T=571640 870360 1 180 $X=567920 $Y=869980
X2659 3280 3262 3324 3336 1 3346 2 AOI22S $T=569160 840120 1 0 $X=569160 $Y=834700
X2660 3210 3202 3335 3019 1 3355 2 AOI22S $T=570400 749400 0 0 $X=570400 $Y=749020
X2661 497 500 3351 503 1 505 2 AOI22S $T=572260 729240 1 0 $X=572260 $Y=723820
X2662 3210 3202 3309 491 1 499 2 AOI22S $T=575980 759480 1 180 $X=572260 $Y=759100
X2663 3035 3262 3356 3364 1 508 2 AOI22S $T=574120 779640 0 0 $X=574120 $Y=779260
X2664 3210 3202 3361 3381 1 3392 2 AOI22S $T=576600 759480 1 0 $X=576600 $Y=754060
X2665 3401 3408 3373 3386 1 2727 2 AOI22S $T=579700 860280 1 0 $X=579700 $Y=854860
X2666 3035 3262 3368 3334 1 2615 2 AOI22S $T=580320 799800 1 0 $X=580320 $Y=794380
X2667 497 500 3416 523 1 528 2 AOI22S $T=582800 739320 0 0 $X=582800 $Y=738940
X2668 3210 494 3372 504 1 526 2 AOI22S $T=582800 779640 1 0 $X=582800 $Y=774220
X2669 532 525 3406 3409 1 2533 2 AOI22S $T=586520 880440 1 180 $X=582800 $Y=880060
X2670 3404 3408 3379 515 1 3402 2 AOI22S $T=584040 840120 1 0 $X=584040 $Y=834700
X2671 3404 494 3431 3438 1 3375 2 AOI22S $T=589000 779640 1 0 $X=589000 $Y=774220
X2672 3401 3408 3424 2321 1 535 2 AOI22S $T=589000 860280 0 0 $X=589000 $Y=859900
X2673 3475 3461 3434 3433 1 2586 2 AOI22S $T=596440 860280 1 180 $X=592720 $Y=859900
X2674 3401 525 3471 3313 1 3456 2 AOI22S $T=595820 880440 1 0 $X=595820 $Y=875020
X2675 3475 3472 3460 2601 1 3492 2 AOI22S $T=597680 840120 1 0 $X=597680 $Y=834700
X2676 3475 3472 3412 3497 1 3449 2 AOI22S $T=598920 819960 0 0 $X=598920 $Y=819580
X2677 3475 3472 3394 3502 1 3342 2 AOI22S $T=599540 830040 0 0 $X=599540 $Y=829660
X2678 3475 3461 3468 549 1 3489 2 AOI22S $T=600160 860280 1 0 $X=600160 $Y=854860
X2679 3475 3461 3369 3517 1 3521 2 AOI22S $T=601400 860280 0 0 $X=601400 $Y=859900
X2680 547 3461 3440 531 1 552 2 AOI22S $T=601400 890520 0 0 $X=601400 $Y=890140
X2681 547 3461 3504 2561 1 3525 2 AOI22S $T=602020 890520 1 0 $X=602020 $Y=885100
X2682 3585 3577 3579 3513 1 3564 2 AOI22S $T=618760 759480 0 180 $X=615040 $Y=754060
X2683 3585 3577 3573 558 1 566 2 AOI22S $T=618760 759480 1 180 $X=615040 $Y=759100
X2684 571 569 3583 568 1 567 2 AOI22S $T=619380 729240 0 180 $X=615660 $Y=723820
X2685 571 569 3594 3469 1 575 2 AOI22S $T=619380 729240 0 0 $X=619380 $Y=728860
X2686 3585 3577 3590 3568 1 3547 2 AOI22S $T=620620 749400 0 0 $X=620620 $Y=749020
X2687 3623 3608 3618 3586 1 574 2 AOI22S $T=624340 779640 0 180 $X=620620 $Y=774220
X2688 3623 3608 3619 3602 1 2751 2 AOI22S $T=624340 779640 1 180 $X=620620 $Y=779260
X2689 3623 3608 3620 3612 1 2642 2 AOI22S $T=625580 789720 0 180 $X=621860 $Y=784300
X2690 3585 3577 3625 584 1 3634 2 AOI22S $T=623720 759480 1 0 $X=623720 $Y=754060
X2691 3637 3628 3631 3500 1 581 2 AOI22S $T=627440 799800 1 180 $X=623720 $Y=799420
X2692 3637 3628 3633 3559 1 595 2 AOI22S $T=628060 799800 1 0 $X=628060 $Y=794380
X2693 571 569 3635 3610 1 585 2 AOI22S $T=628680 729240 0 0 $X=628680 $Y=728860
X2694 3637 3628 3639 614 1 616 2 AOI22S $T=637360 799800 1 0 $X=637360 $Y=794380
X2695 3585 3577 3694 628 1 3670 2 AOI22S $T=642320 759480 1 0 $X=642320 $Y=754060
X2696 3623 3608 3700 3695 1 2662 2 AOI22S $T=645420 779640 1 0 $X=645420 $Y=774220
X2697 3637 3628 3705 3709 1 3651 2 AOI22S $T=646660 799800 0 0 $X=646660 $Y=799420
X2698 635 3746 3740 638 1 632 2 AOI22S $T=650380 729240 1 0 $X=650380 $Y=723820
X2699 3623 3608 3753 3754 1 3727 2 AOI22S $T=655340 779640 0 180 $X=651620 $Y=774220
X2700 3767 3748 3770 3758 1 602 2 AOI22S $T=655340 840120 0 180 $X=651620 $Y=834700
X2701 644 642 3772 3661 1 599 2 AOI22S $T=655340 890520 1 180 $X=651620 $Y=890140
X2702 3767 3748 3775 3675 1 3701 2 AOI22S $T=656580 830040 1 180 $X=652860 $Y=829660
X2703 3773 3628 3747 3682 1 648 2 AOI22S $T=655340 799800 0 0 $X=655340 $Y=799420
X2704 3767 3778 3782 3766 1 3658 2 AOI22S $T=659060 850200 0 180 $X=655340 $Y=844780
X2705 3767 3778 3795 3751 1 621 2 AOI22S $T=660920 870360 0 180 $X=657200 $Y=864940
X2706 3773 3778 3802 3793 1 3689 2 AOI22S $T=662160 880440 0 180 $X=658440 $Y=875020
X2707 3767 3778 3792 3812 1 630 2 AOI22S $T=659060 850200 1 0 $X=659060 $Y=844780
X2708 3767 3778 3813 3588 1 631 2 AOI22S $T=664640 870360 0 180 $X=660920 $Y=864940
X2709 635 3746 3816 658 1 657 2 AOI22S $T=665880 729240 0 180 $X=662160 $Y=723820
X2710 3739 3735 3839 660 1 3819 2 AOI22S $T=669600 749400 1 0 $X=669600 $Y=743980
X2711 3796 3842 3841 3845 1 3854 2 AOI22S $T=669600 769560 1 0 $X=669600 $Y=764140
X2712 635 661 3857 679 1 682 2 AOI22S $T=673320 729240 0 0 $X=673320 $Y=728860
X2713 3739 3735 3862 667 1 3790 2 AOI22S $T=673320 749400 1 0 $X=673320 $Y=743980
X2714 3785 3748 3868 3776 1 3826 2 AOI22S $T=677040 799800 0 180 $X=673320 $Y=794380
X2715 3896 3902 3893 3865 1 3284 2 AOI22S $T=683240 840120 0 180 $X=679520 $Y=834700
X2716 3921 3903 3895 3560 1 3905 2 AOI22S $T=684480 850200 1 180 $X=680760 $Y=849820
X2717 3921 3903 3922 665 1 3703 2 AOI22S $T=685100 870360 0 180 $X=681380 $Y=864940
X2718 3739 3735 3919 694 1 3885 2 AOI22S $T=685720 749400 0 180 $X=682000 $Y=743980
X2719 3921 3903 3926 3849 1 693 2 AOI22S $T=686960 880440 0 180 $X=683240 $Y=875020
X2720 635 661 3918 699 1 700 2 AOI22S $T=685100 729240 0 0 $X=685100 $Y=728860
X2721 3898 3842 3937 3929 1 3860 2 AOI22S $T=688820 769560 1 180 $X=685100 $Y=769180
X2722 3921 3935 3931 3814 1 3932 2 AOI22S $T=685720 870360 1 0 $X=685720 $Y=864940
X2723 3921 3935 3925 3728 1 703 2 AOI22S $T=686340 850200 1 0 $X=686340 $Y=844780
X2724 3785 3888 3936 3953 1 3961 2 AOI22S $T=688820 799800 1 0 $X=688820 $Y=794380
X2725 3896 3902 3954 3876 1 3944 2 AOI22S $T=690060 819960 0 0 $X=690060 $Y=819580
X2726 3739 3735 3958 3963 1 3952 2 AOI22S $T=694400 749400 0 180 $X=690680 $Y=743980
X2727 4035 4014 3964 3985 1 4008 2 AOI22S $T=702460 890520 1 180 $X=698740 $Y=890140
X2728 3999 4012 3847 4019 1 4029 2 AOI22S $T=699360 819960 1 0 $X=699360 $Y=814540
X2729 4016 4012 3873 4044 1 4029 2 AOI22S $T=700600 809880 0 0 $X=700600 $Y=809500
X2730 3785 3888 4051 4037 1 3987 2 AOI22S $T=706800 799800 0 180 $X=703080 $Y=794380
X2731 4031 4012 3846 4042 1 4029 2 AOI22S $T=703080 819960 1 0 $X=703080 $Y=814540
X2732 4041 4054 3872 4012 1 4029 2 AOI22S $T=704940 809880 0 0 $X=704940 $Y=809500
X2733 4027 4039 4065 4015 1 4023 2 AOI22S $T=709280 749400 1 180 $X=705560 $Y=749020
X2734 4035 4014 3988 4068 1 4056 2 AOI22S $T=706180 870360 0 0 $X=706180 $Y=869980
X2735 3785 3888 4066 4082 1 4077 2 AOI22S $T=707420 799800 1 0 $X=707420 $Y=794380
X2736 4069 4012 4061 4098 1 4029 2 AOI22S $T=708660 809880 0 0 $X=708660 $Y=809500
X2737 4033 661 4046 729 1 740 2 AOI22S $T=709900 729240 0 0 $X=709900 $Y=728860
X2738 3898 3842 4081 742 1 4095 2 AOI22S $T=710520 769560 1 0 $X=710520 $Y=764140
X2739 4118 4107 4097 745 1 4089 2 AOI22S $T=717340 830040 1 180 $X=713620 $Y=829660
X2740 4027 4039 4099 4113 1 4122 2 AOI22S $T=714240 749400 0 0 $X=714240 $Y=749020
X2741 4118 4107 4120 4111 1 4091 2 AOI22S $T=717960 819960 0 180 $X=714240 $Y=814540
X2742 4189 4196 4086 4217 1 4227 2 AOI22S $T=735320 819960 0 0 $X=735320 $Y=819580
X2743 4189 4196 4125 4223 1 794 2 AOI22S $T=735940 819960 1 0 $X=735940 $Y=814540
X2744 4189 4196 4071 4228 1 4184 2 AOI22S $T=736560 850200 0 0 $X=736560 $Y=849820
X2745 790 793 4004 4247 1 4249 2 AOI22S $T=740280 880440 1 0 $X=740280 $Y=875020
X2746 790 793 4100 807 1 4248 2 AOI22S $T=741520 870360 1 0 $X=741520 $Y=864940
X2747 861 4394 4397 4325 1 4369 2 AOI22S $T=772520 850200 1 180 $X=768800 $Y=849820
X2748 861 857 4415 4358 1 4343 2 AOI22S $T=773140 890520 0 180 $X=769420 $Y=885100
X2749 4400 4412 4429 845 1 852 2 AOI22S $T=776860 799800 1 180 $X=773140 $Y=799420
X2750 861 857 4430 866 1 4392 2 AOI22S $T=776860 890520 1 180 $X=773140 $Y=890140
X2751 4402 4399 4440 4447 1 4416 2 AOI22S $T=776240 759480 1 0 $X=776240 $Y=754060
X2752 861 4394 4446 4258 1 4341 2 AOI22S $T=776860 860280 0 0 $X=776860 $Y=859900
X2753 4400 4412 4464 844 1 4443 2 AOI22S $T=783680 809880 0 180 $X=779960 $Y=804460
X2754 4400 4412 4473 4470 1 882 2 AOI22S $T=786160 819960 0 180 $X=782440 $Y=814540
X2755 4427 4399 4492 864 1 870 2 AOI22S $T=787400 759480 0 180 $X=783680 $Y=754060
X2756 4474 4485 4477 886 1 4468 2 AOI22S $T=783680 840120 1 0 $X=783680 $Y=834700
X2757 4495 4485 4500 4510 1 4513 2 AOI22S $T=787400 799800 0 0 $X=787400 $Y=799420
X2758 4474 897 4524 4453 1 4482 2 AOI22S $T=792360 890520 0 180 $X=788640 $Y=885100
X2759 4379 4396 4514 884 1 894 2 AOI22S $T=791120 749400 1 0 $X=791120 $Y=743980
X2760 4540 897 4546 896 1 898 2 AOI22S $T=794840 860280 1 180 $X=791120 $Y=859900
X2761 4427 4399 4527 902 1 4511 2 AOI22S $T=792360 759480 0 0 $X=792360 $Y=759100
X2762 4379 4396 4532 4486 1 4574 2 AOI22S $T=794840 749400 1 0 $X=794840 $Y=743980
X2763 4495 4485 4535 4335 1 4362 2 AOI22S $T=796700 799800 1 0 $X=796700 $Y=794380
X2764 4474 897 4593 918 1 919 2 AOI22S $T=801660 890520 0 0 $X=801660 $Y=890140
X2765 4379 4396 4497 4588 1 920 2 AOI22S $T=802280 749400 0 0 $X=802280 $Y=749020
X2766 4495 4485 4603 4501 1 914 2 AOI22S $T=802900 819960 0 0 $X=802900 $Y=819580
X2767 4700 4396 4677 4723 1 935 2 AOI22S $T=819640 759480 1 0 $X=819640 $Y=754060
X2768 4427 4721 4713 4567 1 4670 2 AOI22S $T=822120 840120 1 0 $X=822120 $Y=834700
X2769 4739 4628 4754 4629 1 4691 2 AOI22S $T=830180 799800 0 180 $X=826460 $Y=794380
X2770 4736 951 4748 946 1 4730 2 AOI22S $T=828320 860280 1 0 $X=828320 $Y=854860
X2771 4736 951 4753 4705 1 4737 2 AOI22S $T=829560 870360 1 0 $X=829560 $Y=864940
X2772 4666 4394 4760 4554 1 4565 2 AOI22S $T=830800 809880 1 0 $X=830800 $Y=804460
X2773 4720 4721 4783 4779 1 4744 2 AOI22S $T=833280 759480 0 0 $X=833280 $Y=759100
X2774 4720 4791 4772 4735 1 4522 2 AOI22S $T=833280 840120 1 0 $X=833280 $Y=834700
X2775 4736 951 4782 4749 1 4798 2 AOI22S $T=833900 890520 0 0 $X=833900 $Y=890140
X2776 4736 951 4758 4763 1 4531 2 AOI22S $T=834520 890520 1 0 $X=834520 $Y=885100
X2777 4824 4800 4701 4812 1 4611 2 AOI22S $T=841960 840120 0 180 $X=838240 $Y=834700
X2778 967 966 4752 4825 1 4598 2 AOI22S $T=843820 880440 1 180 $X=840100 $Y=880060
X2779 967 966 4773 4831 1 4835 2 AOI22S $T=841340 890520 0 0 $X=841340 $Y=890140
X2780 4739 4802 4826 4836 1 4842 2 AOI22S $T=842580 799800 1 0 $X=842580 $Y=794380
X2781 4824 966 4743 969 1 4313 2 AOI22S $T=843200 880440 1 0 $X=843200 $Y=875020
X2782 4824 966 4746 4472 1 4719 2 AOI22S $T=844440 860280 0 0 $X=844440 $Y=859900
X2783 4700 4849 4854 4817 1 4818 2 AOI22S $T=848780 739320 1 180 $X=845060 $Y=738940
X2784 4720 4721 4859 4848 1 4808 2 AOI22S $T=849400 759480 1 180 $X=845680 $Y=759100
X2785 4890 4849 4867 970 1 4768 2 AOI22S $T=851880 739320 0 180 $X=848160 $Y=733900
X2786 4666 4863 4856 4805 1 4858 2 AOI22S $T=848160 819960 1 0 $X=848160 $Y=814540
X2787 4908 4893 4879 4934 1 4922 2 AOI22S $T=858080 749400 0 0 $X=858080 $Y=749020
X2788 4915 4912 4929 4757 1 4671 2 AOI22S $T=862420 840120 0 180 $X=858700 $Y=834700
X2789 4908 4893 4955 984 1 4898 2 AOI22S $T=866140 749400 1 180 $X=862420 $Y=749020
X2790 4739 4802 4950 4943 1 4926 2 AOI22S $T=867380 789720 0 180 $X=863660 $Y=784300
X2791 4968 4802 4961 4956 1 4875 2 AOI22S $T=869860 809880 0 180 $X=866140 $Y=804460
X2792 4739 4802 4965 4958 1 4637 2 AOI22S $T=870480 789720 1 180 $X=866760 $Y=789340
X2793 4890 4918 4957 4959 1 989 2 AOI22S $T=871100 729240 1 180 $X=867380 $Y=728860
X2794 4982 4981 4977 4942 1 4907 2 AOI22S $T=873580 850200 1 180 $X=869860 $Y=849820
X2795 4908 4893 5038 5004 1 4994 2 AOI22S $T=880400 749400 1 180 $X=876680 $Y=749020
X2796 4890 4918 5041 1002 1 5015 2 AOI22S $T=882260 739320 0 180 $X=878540 $Y=733900
X2797 4915 4912 5049 5046 1 5083 2 AOI22S $T=883500 850200 0 0 $X=883500 $Y=849820
X2798 4908 4893 5070 1007 1 4983 2 AOI22S $T=887840 749400 1 180 $X=884120 $Y=749020
X2799 4908 4893 5081 5087 1 5069 2 AOI22S $T=887840 749400 0 0 $X=887840 $Y=749020
X2800 4890 4918 5103 1021 1 1013 2 AOI22S $T=892800 739320 1 0 $X=892800 $Y=733900
X2801 4982 4981 5073 5132 1 5121 2 AOI22S $T=896520 860280 1 0 $X=896520 $Y=854860
X2802 4982 4981 5089 5142 1 5170 2 AOI22S $T=897760 880440 1 0 $X=897760 $Y=875020
X2803 4982 4981 5017 5147 1 5157 2 AOI22S $T=899000 870360 0 0 $X=899000 $Y=869980
X2804 4982 4981 5062 5166 1 5144 2 AOI22S $T=900240 860280 1 0 $X=900240 $Y=854860
X2805 5295 5287 5289 5235 1 5275 2 AOI22S $T=930620 769560 1 180 $X=926900 $Y=769180
X2806 5326 5309 5308 5241 1 5268 2 AOI22S $T=933720 759480 0 180 $X=930000 $Y=754060
X2807 5319 5307 5303 5301 1 5299 2 AOI22S $T=933720 830040 0 180 $X=930000 $Y=824620
X2808 5328 5316 5311 5237 1 5283 2 AOI22S $T=934960 799800 0 180 $X=931240 $Y=794380
X2809 5332 5324 5363 1047 1 5305 2 AOI22S $T=936820 880440 1 180 $X=933100 $Y=880060
X2810 5326 5355 5375 5342 1 5310 2 AOI22S $T=941160 759480 0 180 $X=937440 $Y=754060
X2811 1067 5356 5369 5360 1 5350 2 AOI22S $T=942400 860280 0 180 $X=938680 $Y=854860
X2812 5328 5316 5362 5321 1 5372 2 AOI22S $T=939300 799800 1 0 $X=939300 $Y=794380
X2813 5295 5287 5364 1061 1 5371 2 AOI22S $T=939920 739320 0 0 $X=939920 $Y=738940
X2814 1051 5293 5394 5348 1 5366 2 AOI22S $T=946120 850200 0 180 $X=942400 $Y=844780
X2815 5257 5385 5370 5358 1 5377 2 AOI22S $T=947360 779640 1 180 $X=943640 $Y=779260
X2816 5332 5324 5415 5400 1 5401 2 AOI22S $T=947360 870360 0 0 $X=947360 $Y=869980
X2817 5326 5316 5420 5396 1 1072 2 AOI22S $T=948600 789720 0 0 $X=948600 $Y=789340
X2818 5445 5307 5417 5329 1 5347 2 AOI22S $T=953560 830040 0 180 $X=949840 $Y=824620
X2819 5437 5356 5438 5410 1 5457 2 AOI22S $T=952320 850200 1 0 $X=952320 $Y=844780
X2820 5319 5385 5422 5481 1 5453 2 AOI22S $T=953560 779640 0 0 $X=953560 $Y=779260
X2821 1078 5468 5412 5472 1 5479 2 AOI22S $T=955420 870360 0 0 $X=955420 $Y=869980
X2822 5332 5324 5473 5482 1 5483 2 AOI22S $T=956660 880440 1 0 $X=956660 $Y=875020
X2823 5461 5287 5484 1084 1 5474 2 AOI22S $T=961000 739320 0 180 $X=957280 $Y=733900
X2824 5319 5385 5488 5444 1 5469 2 AOI22S $T=961620 779640 1 180 $X=957900 $Y=779260
X2825 5319 5385 5515 5530 1 5532 2 AOI22S $T=965340 779640 0 0 $X=965340 $Y=779260
X2826 5332 5468 5512 5535 1 5540 2 AOI22S $T=966580 880440 1 0 $X=966580 $Y=875020
X2827 5328 5316 5537 5513 1 5551 2 AOI22S $T=968440 799800 1 0 $X=968440 $Y=794380
X2828 5437 5356 5523 5465 1 5547 2 AOI22S $T=968440 840120 0 0 $X=968440 $Y=839740
X2829 1051 1093 5538 5543 1 1095 2 AOI22S $T=968440 890520 1 0 $X=968440 $Y=885100
X2830 5437 5356 5565 5607 1 5579 2 AOI22S $T=972780 840120 0 0 $X=972780 $Y=839740
X2831 1078 5468 5548 5573 1 5582 2 AOI22S $T=972780 880440 1 0 $X=972780 $Y=875020
X2832 5475 5355 5563 5518 1 5598 2 AOI22S $T=975260 759480 1 0 $X=975260 $Y=754060
X2833 5445 5307 5589 5599 1 5603 2 AOI22S $T=975880 830040 0 0 $X=975880 $Y=829660
X2834 5461 5528 5601 5606 1 5612 2 AOI22S $T=977740 739320 0 0 $X=977740 $Y=738940
X2835 5649 5675 5685 5673 1 5647 2 AOI22S $T=999440 809880 0 180 $X=995720 $Y=804460
X2836 1119 5687 5690 5658 1 5679 2 AOI22S $T=1000680 860280 0 180 $X=996960 $Y=854860
X2837 5663 5674 5705 5682 1 5652 2 AOI22S $T=1001300 779640 1 180 $X=997580 $Y=779260
X2838 5689 5716 5717 5656 1 1121 2 AOI22S $T=1004400 739320 1 180 $X=1000680 $Y=738940
X2839 1119 5687 5708 5719 1 1111 2 AOI22S $T=1000680 860280 0 0 $X=1000680 $Y=859900
X2840 5649 5687 5723 5741 1 5737 2 AOI22S $T=1002540 840120 1 0 $X=1002540 $Y=834700
X2841 5649 5675 5730 1127 1 5744 2 AOI22S $T=1003160 799800 0 0 $X=1003160 $Y=799420
X2842 1133 1129 5739 5662 1 5660 2 AOI22S $T=1007500 890520 1 180 $X=1003780 $Y=890140
X2843 1133 5749 5715 1128 1 5641 2 AOI22S $T=1008120 880440 1 180 $X=1004400 $Y=880060
X2844 5689 5749 5761 5645 1 5757 2 AOI22S $T=1009980 880440 0 180 $X=1006260 $Y=875020
X2845 5779 5681 5726 5768 1 5650 2 AOI22S $T=1011840 769560 0 180 $X=1008120 $Y=764140
X2846 5663 5674 5758 5693 1 5784 2 AOI22S $T=1009980 779640 0 0 $X=1009980 $Y=779260
X2847 5778 5716 5748 5777 1 1142 2 AOI22S $T=1011220 739320 0 0 $X=1011220 $Y=738940
X2848 5779 5681 5742 5789 1 5692 2 AOI22S $T=1011840 769560 0 0 $X=1011840 $Y=769180
X2849 5840 5749 5832 5790 1 1139 2 AOI22S $T=1024240 890520 1 180 $X=1020520 $Y=890140
X2850 5845 5675 5838 5835 1 5756 2 AOI22S $T=1024860 850200 0 180 $X=1021140 $Y=844780
X2851 5689 5749 5831 5786 1 5680 2 AOI22S $T=1021760 880440 1 0 $X=1021760 $Y=875020
X2852 5778 5716 5852 5846 1 1155 2 AOI22S $T=1026720 739320 1 180 $X=1023000 $Y=738940
X2853 5779 5681 5861 5812 1 5841 2 AOI22S $T=1027340 769560 0 180 $X=1023620 $Y=764140
X2854 5864 5674 5850 5847 1 5848 2 AOI22S $T=1027960 789720 0 180 $X=1024240 $Y=784300
X2855 5839 5855 5842 5854 1 5844 2 AOI22S $T=1024240 809880 1 0 $X=1024240 $Y=804460
X2856 5845 5687 5851 5806 1 5821 2 AOI22S $T=1024860 860280 1 0 $X=1024860 $Y=854860
X2857 5873 5876 5747 1161 1 1165 2 AOI22S $T=1028580 890520 0 0 $X=1028580 $Y=890140
X2858 5873 5876 5828 1167 1 1163 2 AOI22S $T=1028580 900600 1 0 $X=1028580 $Y=895180
X2859 5839 5855 5896 5882 1 5859 2 AOI22S $T=1033540 809880 1 180 $X=1029820 $Y=809500
X2860 5778 5716 5885 5911 1 1173 2 AOI22S $T=1032920 739320 0 0 $X=1032920 $Y=738940
X2861 5873 5876 5866 5884 1 5920 2 AOI22S $T=1033540 880440 1 0 $X=1033540 $Y=875020
X2862 5873 5876 5709 5914 1 5929 2 AOI22S $T=1034160 890520 1 0 $X=1034160 $Y=885100
X2863 5779 5924 5880 5897 1 5909 2 AOI22S $T=1038500 769560 0 180 $X=1034780 $Y=764140
X2864 5864 5674 5895 5907 1 5933 2 AOI22S $T=1034780 779640 0 0 $X=1034780 $Y=779260
X2865 5941 5876 5767 5925 1 5921 2 AOI22S $T=1039120 850200 1 180 $X=1035400 $Y=849820
X2866 5778 5946 5953 5944 1 1178 2 AOI22S $T=1042840 739320 1 180 $X=1039120 $Y=738940
X2867 5970 5924 5948 5931 1 1182 2 AOI22S $T=1045320 759480 0 180 $X=1041600 $Y=754060
X2868 5845 5675 5954 5962 1 5967 2 AOI22S $T=1041600 850200 1 0 $X=1041600 $Y=844780
X2869 5839 5855 5959 5960 1 5952 2 AOI22S $T=1042220 799800 0 0 $X=1042220 $Y=799420
X2870 5864 5674 5958 5975 1 5936 2 AOI22S $T=1045320 779640 0 0 $X=1045320 $Y=779260
X2871 5970 5924 5987 5986 1 6006 2 AOI22S $T=1048420 759480 0 0 $X=1048420 $Y=759100
X2872 5941 5998 5980 5979 1 5957 2 AOI22S $T=1049040 860280 1 0 $X=1049040 $Y=854860
X2873 5839 5855 6000 6011 1 5990 2 AOI22S $T=1050900 809880 1 0 $X=1050900 $Y=804460
X2874 5840 5704 5982 5981 1 6016 2 AOI22S $T=1050900 880440 1 0 $X=1050900 $Y=875020
X2875 5864 6050 5994 6028 1 6056 2 AOI22S $T=1058340 769560 0 0 $X=1058340 $Y=769180
X2876 5970 5924 6045 6032 1 6067 2 AOI22S $T=1061440 759480 1 0 $X=1061440 $Y=754060
X2877 5864 6050 6053 6054 1 6075 2 AOI22S $T=1062060 769560 0 0 $X=1062060 $Y=769180
X2878 6064 6072 6046 1197 1 1196 2 AOI22S $T=1063920 729240 0 0 $X=1063920 $Y=728860
X2879 1198 1193 6077 6008 1 6055 2 AOI22S $T=1068880 890520 1 180 $X=1065160 $Y=890140
X2880 5941 5998 6068 6062 1 5984 2 AOI22S $T=1070120 860280 0 180 $X=1066400 $Y=854860
X2881 6108 6100 6079 6078 1 6037 2 AOI22S $T=1071360 830040 1 180 $X=1067640 $Y=829660
X2882 6109 5704 6071 6015 1 6094 2 AOI22S $T=1071360 870360 1 180 $X=1067640 $Y=869980
X2883 6099 6136 6138 6129 1 6125 2 AOI22S $T=1079420 809880 0 180 $X=1075700 $Y=804460
X2884 6064 6072 6145 1214 1 1212 2 AOI22S $T=1080660 729240 1 180 $X=1076940 $Y=728860
X2885 5970 5924 6149 6120 1 6139 2 AOI22S $T=1081280 759480 1 180 $X=1077560 $Y=759100
X2886 5941 5998 6151 6133 1 1222 2 AOI22S $T=1080040 860280 1 0 $X=1080040 $Y=854860
X2887 6109 6162 6169 6156 1 6135 2 AOI22S $T=1083760 870360 0 180 $X=1080040 $Y=864940
X2888 6194 6069 6161 6164 1 6092 2 AOI22S $T=1085000 779640 0 180 $X=1081280 $Y=774220
X2889 6108 6100 6183 6085 1 6165 2 AOI22S $T=1085000 830040 0 180 $X=1081280 $Y=824620
X2890 6099 6136 6176 6160 1 6103 2 AOI22S $T=1086240 809880 0 180 $X=1082520 $Y=804460
X2891 6194 6069 6190 6157 1 6174 2 AOI22S $T=1088100 779640 1 0 $X=1088100 $Y=774220
X2892 6109 6162 6201 6223 1 6211 2 AOI22S $T=1089340 870360 1 0 $X=1089340 $Y=864940
X2893 6064 6072 6184 1221 1 1223 2 AOI22S $T=1090580 729240 1 0 $X=1090580 $Y=723820
X2894 6108 6100 6239 6246 1 6238 2 AOI22S $T=1096160 830040 1 0 $X=1096160 $Y=824620
X2895 6194 6069 6242 6232 1 6250 2 AOI22S $T=1096780 779640 1 0 $X=1096780 $Y=774220
X2896 6248 6178 6260 6227 1 6225 2 AOI22S $T=1101740 749400 1 180 $X=1098020 $Y=749020
X2897 6147 5998 6234 6256 1 6263 2 AOI22S $T=1098020 850200 0 0 $X=1098020 $Y=849820
X2898 6064 6072 6235 6259 1 1235 2 AOI22S $T=1098640 729240 1 0 $X=1098640 $Y=723820
X2899 6108 6100 6255 6269 1 6267 2 AOI22S $T=1099260 840120 1 0 $X=1099260 $Y=834700
X2900 6099 6136 6287 6340 1 6297 2 AOI22S $T=1104840 809880 1 0 $X=1104840 $Y=804460
X2901 6064 6072 6311 6310 1 1242 2 AOI22S $T=1111660 739320 0 180 $X=1107940 $Y=733900
X2902 6248 6178 6304 6319 1 6322 2 AOI22S $T=1107940 749400 1 0 $X=1107940 $Y=743980
X2903 6147 1244 6281 6328 1 6329 2 AOI22S $T=1109180 870360 0 0 $X=1109180 $Y=869980
X2904 6109 1236 6286 6323 1 1246 2 AOI22S $T=1109180 880440 1 0 $X=1109180 $Y=875020
X2905 6064 6072 6312 6339 1 1250 2 AOI22S $T=1110420 729240 0 0 $X=1110420 $Y=728860
X2906 3740 3736 3747 3753 2 1 3769 AN4S $T=649760 759480 1 0 $X=649760 $Y=754060
X2907 3816 3839 3844 3841 2 1 3870 AN4S $T=669600 759480 0 0 $X=669600 $Y=759100
X2908 3857 3862 3868 3833 2 1 3880 AN4S $T=673320 749400 0 0 $X=673320 $Y=749020
X2909 3918 3919 3936 3937 2 1 3904 AN4S $T=685720 749400 0 0 $X=685720 $Y=749020
X2910 709 3959 704 3891 2 1 3933 AN4S $T=692540 900600 0 180 $X=687580 $Y=895180
X2911 3966 3964 3772 3907 2 1 3942 AN4S $T=693160 890520 1 180 $X=688200 $Y=890140
X2912 705 3958 3965 3969 2 1 3960 AN4S $T=690680 759480 0 0 $X=690680 $Y=759100
X2913 4004 3995 3802 3926 2 1 3979 AN4S $T=699360 880440 0 180 $X=694400 $Y=875020
X2914 3988 3931 3795 4003 2 1 4002 AN4S $T=696260 870360 1 0 $X=696260 $Y=864940
X2915 4065 4052 4051 4046 2 1 3982 AN4S $T=708660 759480 0 180 $X=703700 $Y=754060
X2916 4093 4099 4066 4081 2 1 4040 AN4S $T=714860 759480 1 180 $X=709900 $Y=759100
X2917 5024 5025 5018 4950 2 1 4963 AN4S $T=881020 789720 1 180 $X=876060 $Y=789340
X2918 5036 5037 5044 1011 2 1 5080 AN4S $T=881020 890520 1 0 $X=881020 $Y=885100
X2919 5102 5091 5086 4965 2 1 5052 AN4S $T=891560 789720 1 180 $X=886600 $Y=789340
X2920 5106 5112 5119 4964 2 1 5129 AN4S $T=893420 789720 1 0 $X=893420 $Y=784300
X2921 5130 5141 5131 4961 2 1 5111 AN4S $T=900860 809880 0 180 $X=895900 $Y=804460
X2922 5151 5154 5159 4974 2 1 5172 AN4S $T=900860 809880 1 0 $X=900860 $Y=804460
X2923 5708 1124 5715 5709 2 1 5359 AN4S $T=1004400 880440 1 180 $X=999440 $Y=880060
X2924 5685 5705 5717 5726 2 1 5569 AN4S $T=1000680 779640 1 0 $X=1000680 $Y=774220
X2925 5690 1125 5739 5747 2 1 5527 AN4S $T=1003160 900600 1 0 $X=1003160 $Y=895180
X2926 5730 5758 5748 5742 2 1 5378 AN4S $T=1008740 779640 1 180 $X=1003780 $Y=779260
X2927 5723 1132 5761 5767 2 1 5424 AN4S $T=1006260 860280 0 0 $X=1006260 $Y=859900
X2928 5838 1156 5832 5828 2 1 1086 AN4S $T=1024860 900600 0 180 $X=1019900 $Y=895180
X2929 5842 5850 5852 5861 2 1 5406 AN4S $T=1024860 779640 0 0 $X=1024860 $Y=779260
X2930 5851 1160 5831 5866 2 1 5373 AN4S $T=1030440 880440 0 180 $X=1025480 $Y=875020
X2931 5896 5895 5885 5880 2 1 5333 AN4S $T=1033540 769560 0 180 $X=1028580 $Y=764140
X2932 5959 5958 5953 5948 2 1 5554 AN4S $T=1044080 779640 1 180 $X=1039120 $Y=779260
X2933 5954 1188 5982 5980 2 1 5428 AN4S $T=1049040 860280 0 180 $X=1044080 $Y=854860
X2934 6000 5994 5988 5987 2 1 5621 AN4S $T=1050900 769560 0 180 $X=1045940 $Y=764140
X2935 6060 6053 6046 6045 2 1 5575 AN4S $T=1061440 759480 1 180 $X=1056480 $Y=759100
X2936 6079 6077 6071 6068 2 1 5320 AN4S $T=1066400 860280 1 180 $X=1061440 $Y=859900
X2937 6138 6161 6145 6149 2 1 5382 AN4S $T=1083140 769560 0 180 $X=1078180 $Y=764140
X2938 6183 6187 6169 6151 2 1 5458 AN4S $T=1088720 860280 0 180 $X=1083760 $Y=854860
X2939 6176 6190 6184 6179 2 1 5318 AN4S $T=1089340 749400 1 180 $X=1084380 $Y=749020
X2940 6209 6216 6202 6199 2 1 5511 AN4S $T=1093680 860280 0 180 $X=1088720 $Y=854860
X2941 6243 6242 6235 6231 2 1 5499 AN4S $T=1098640 759480 0 180 $X=1093680 $Y=754060
X2942 6239 1231 6201 6234 2 1 5605 AN4S $T=1098640 860280 0 180 $X=1093680 $Y=854860
X2943 6275 1239 6285 6281 2 1 5558 AN4S $T=1107940 870360 1 180 $X=1102980 $Y=869980
X2944 6255 1240 6286 6282 2 1 5418 AN4S $T=1107940 880440 1 180 $X=1102980 $Y=880060
X2945 6287 6306 6311 6260 2 1 5421 AN4S $T=1111660 759480 0 180 $X=1106700 $Y=754060
X2946 6284 6305 6312 6304 2 1 5594 AN4S $T=1107320 759480 0 0 $X=1107320 $Y=759100
X2947 1418 2 1 1412 BUF1 $T=234980 779640 0 0 $X=234980 $Y=779260
X2948 51 2 1 58 BUF1 $T=254200 739320 1 0 $X=254200 $Y=733900
X2949 1547 2 1 1396 BUF1 $T=262260 789720 0 180 $X=259780 $Y=784300
X2950 1650 2 1 1433 BUF1 $T=280240 799800 0 180 $X=277760 $Y=794380
X2951 76 2 1 98 BUF1 $T=285200 819960 1 0 $X=285200 $Y=814540
X2952 97 2 1 1677 BUF1 $T=287060 729240 0 0 $X=287060 $Y=728860
X2953 78 2 1 113 BUF1 $T=295120 819960 1 0 $X=295120 $Y=814540
X2954 120 2 1 1714 BUF1 $T=305040 830040 0 180 $X=302560 $Y=824620
X2955 120 2 1 1878 BUF1 $T=314960 830040 1 0 $X=314960 $Y=824620
X2956 163 2 1 138 BUF1 $T=322400 729240 0 180 $X=319920 $Y=723820
X2957 120 2 1 163 BUF1 $T=326120 729240 0 180 $X=323640 $Y=723820
X2958 120 2 1 1970 BUF1 $T=329220 830040 1 0 $X=329220 $Y=824620
X2959 158 2 1 2153 BUF1 $T=361460 840120 0 0 $X=361460 $Y=839740
X2960 2067 2 1 2194 BUF1 $T=362700 789720 0 0 $X=362700 $Y=789340
X2961 1871 2 1 2189 BUF1 $T=367660 840120 1 0 $X=367660 $Y=834700
X2962 235 2 1 2390 BUF1 $T=394320 830040 1 0 $X=394320 $Y=824620
X2963 269 2 1 2603 BUF1 $T=430900 870360 1 0 $X=430900 $Y=864940
X2964 2305 2 1 2641 BUF1 $T=442680 799800 1 0 $X=442680 $Y=794380
X2965 2155 2 1 338 BUF1 $T=445160 819960 1 180 $X=442680 $Y=819580
X2966 2641 2 1 337 BUF1 $T=447020 870360 1 0 $X=447020 $Y=864940
X2967 2706 2 1 345 BUF1 $T=451980 860280 0 180 $X=449500 $Y=854860
X2968 2739 2 1 2674 BUF1 $T=458180 799800 1 0 $X=458180 $Y=794380
X2969 2786 2 1 2699 BUF1 $T=466860 779640 1 180 $X=464380 $Y=779260
X2970 2824 2 1 366 BUF1 $T=475540 880440 1 180 $X=473060 $Y=880060
X2971 2756 2 1 2700 BUF1 $T=476160 840120 1 0 $X=476160 $Y=834700
X2972 2879 2 1 2689 BUF1 $T=487940 799800 0 180 $X=485460 $Y=794380
X2973 2895 2 1 2756 BUF1 $T=489180 850200 1 0 $X=489180 $Y=844780
X2974 2929 2 1 2739 BUF1 $T=496000 799800 0 0 $X=496000 $Y=799420
X2975 2155 2 1 409 BUF1 $T=498480 749400 1 0 $X=498480 $Y=743980
X2976 2993 2 1 2786 BUF1 $T=502200 789720 1 180 $X=499720 $Y=789340
X2977 411 2 1 2857 BUF1 $T=503440 809880 0 180 $X=500960 $Y=804460
X2978 420 2 1 2929 BUF1 $T=505920 900600 1 0 $X=505920 $Y=895180
X2979 3021 2 1 2843 BUF1 $T=512740 840120 0 180 $X=510260 $Y=834700
X2980 3045 2 1 2931 BUF1 $T=518320 769560 0 180 $X=515840 $Y=764140
X2981 433 2 1 2824 BUF1 $T=518320 870360 0 180 $X=515840 $Y=864940
X2982 3077 2 1 2879 BUF1 $T=525760 799800 1 180 $X=523280 $Y=799420
X2983 3077 2 1 423 BUF1 $T=526380 890520 0 0 $X=526380 $Y=890140
X2984 3137 2 1 433 BUF1 $T=531960 789720 0 180 $X=529480 $Y=784300
X2985 3202 2 1 3084 BUF1 $T=546220 759480 0 180 $X=543740 $Y=754060
X2986 2963 2 1 3211 BUF1 $T=546220 729240 0 0 $X=546220 $Y=728860
X2987 3210 2 1 3099 BUF1 $T=549320 749400 1 180 $X=546840 $Y=749020
X2988 2831 2 1 3233 BUF1 $T=549320 749400 1 0 $X=549320 $Y=743980
X2989 3211 2 1 459 BUF1 $T=557380 729240 0 180 $X=554900 $Y=723820
X2990 3151 2 1 3263 BUF1 $T=561100 779640 0 0 $X=561100 $Y=779260
X2991 482 2 1 3297 BUF1 $T=561720 890520 1 0 $X=561720 $Y=885100
X2992 495 2 1 1969 BUF1 $T=571020 819960 0 180 $X=568540 $Y=814540
X2993 3297 2 1 3262 BUF1 $T=571020 840120 1 180 $X=568540 $Y=839740
X2994 3015 2 1 3352 BUF1 $T=571020 840120 0 0 $X=571020 $Y=839740
X2995 3401 2 1 532 BUF1 $T=586520 880440 0 0 $X=586520 $Y=880060
X2996 3404 2 1 3401 BUF1 $T=589620 850200 1 0 $X=589620 $Y=844780
X2997 2987 2 1 537 BUF1 $T=590240 749400 1 0 $X=590240 $Y=743980
X2998 541 2 1 2260 BUF1 $T=593960 779640 0 0 $X=593960 $Y=779260
X2999 3225 2 1 3250 BUF1 $T=593960 799800 0 0 $X=593960 $Y=799420
X3000 3472 2 1 544 BUF1 $T=595820 900600 1 0 $X=595820 $Y=895180
X3001 3015 2 1 3487 BUF1 $T=597060 799800 0 0 $X=597060 $Y=799420
X3002 3225 2 1 529 BUF1 $T=600160 739320 0 0 $X=600160 $Y=738940
X3003 3186 2 1 3593 BUF1 $T=617520 890520 1 0 $X=617520 $Y=885100
X3004 3316 2 1 3609 BUF1 $T=623720 840120 1 0 $X=623720 $Y=834700
X3005 3482 2 1 591 BUF1 $T=625580 850200 1 0 $X=625580 $Y=844780
X3006 560 2 1 3652 BUF1 $T=642940 779640 1 0 $X=642940 $Y=774220
X3007 3739 2 1 3585 BUF1 $T=649140 749400 1 180 $X=646660 $Y=749020
X3008 3748 2 1 3628 BUF1 $T=652860 799800 1 180 $X=650380 $Y=799420
X3009 3761 2 1 3773 BUF1 $T=652860 799800 0 0 $X=652860 $Y=799420
X3010 3778 2 1 3748 BUF1 $T=658440 840120 1 180 $X=655960 $Y=839740
X3011 3791 2 1 3486 BUF1 $T=660920 779640 1 180 $X=658440 $Y=779260
X3012 3796 2 1 3623 BUF1 $T=661540 769560 0 180 $X=659060 $Y=764140
X3013 642 2 1 3778 BUF1 $T=659060 890520 0 0 $X=659060 $Y=890140
X3014 661 2 1 3746 BUF1 $T=668360 729240 0 180 $X=665880 $Y=723820
X3015 3652 2 1 676 BUF1 $T=670220 850200 1 0 $X=670220 $Y=844780
X3016 428 2 1 677 BUF1 $T=672700 729240 1 0 $X=672700 $Y=723820
X3017 3511 2 1 681 BUF1 $T=672700 890520 0 0 $X=672700 $Y=890140
X3018 3898 2 1 3796 BUF1 $T=682000 769560 1 180 $X=679520 $Y=769180
X3019 3902 2 1 3903 BUF1 $T=684480 830040 1 180 $X=682000 $Y=829660
X3020 426 2 1 3875 BUF1 $T=687580 759480 0 0 $X=687580 $Y=759100
X3021 3994 2 1 654 BUF1 $T=699360 819960 1 180 $X=696880 $Y=819580
X3022 3593 2 1 728 BUF1 $T=700600 880440 1 0 $X=700600 $Y=875020
X3023 4033 2 1 635 BUF1 $T=704320 729240 0 180 $X=701840 $Y=723820
X3024 3902 2 1 3842 BUF1 $T=704320 769560 1 180 $X=701840 $Y=769180
X3025 4014 2 1 730 BUF1 $T=703700 890520 0 0 $X=703700 $Y=890140
X3026 4035 2 1 731 BUF1 $T=704320 900600 1 0 $X=704320 $Y=895180
X3027 3233 2 1 732 BUF1 $T=708660 729240 1 0 $X=708660 $Y=723820
X3028 4107 2 1 4039 BUF1 $T=716720 769560 0 180 $X=714240 $Y=764140
X3029 4107 2 1 4014 BUF1 $T=714240 840120 0 0 $X=714240 $Y=839740
X3030 625 2 1 752 BUF1 $T=714860 900600 1 0 $X=714860 $Y=895180
X3031 4118 2 1 4035 BUF1 $T=715480 850200 1 0 $X=715480 $Y=844780
X3032 4189 2 1 4033 BUF1 $T=734080 779640 0 180 $X=731600 $Y=774220
X3033 4196 2 1 661 BUF1 $T=736560 769560 1 180 $X=734080 $Y=769180
X3034 4244 2 1 253 BUF1 $T=740280 799800 0 0 $X=740280 $Y=799420
X3035 4189 2 1 790 BUF1 $T=744000 850200 1 180 $X=741520 $Y=849820
X3036 4196 2 1 793 BUF1 $T=745240 860280 0 180 $X=742760 $Y=854860
X3037 813 2 1 3165 BUF1 $T=747100 799800 1 180 $X=744620 $Y=799420
X3038 819 2 1 815 BUF1 $T=748960 799800 0 180 $X=746480 $Y=794380
X3039 4178 2 1 4357 BUF1 $T=766940 860280 0 180 $X=764460 $Y=854860
X3040 4384 2 1 4252 BUF1 $T=770040 769560 1 180 $X=767560 $Y=769180
X3041 857 2 1 4394 BUF1 $T=768800 809880 1 0 $X=768800 $Y=804460
X3042 3859 2 1 4370 BUF1 $T=770040 860280 0 0 $X=770040 $Y=859900
X3043 4402 2 1 4427 BUF1 $T=773760 759480 1 0 $X=773760 $Y=754060
X3044 4243 2 1 4437 BUF1 $T=773760 830040 0 0 $X=773760 $Y=829660
X3045 867 2 1 4047 BUF1 $T=775000 779640 1 0 $X=775000 $Y=774220
X3046 4144 2 1 4454 BUF1 $T=777480 809880 1 0 $X=777480 $Y=804460
X3047 4338 2 1 4434 BUF1 $T=780580 779640 0 0 $X=780580 $Y=779260
X3048 4437 2 1 881 BUF1 $T=781820 799800 0 0 $X=781820 $Y=799420
X3049 4370 2 1 4480 BUF1 $T=781820 860280 0 0 $X=781820 $Y=859900
X3050 4485 2 1 897 BUF1 $T=788640 860280 0 0 $X=788640 $Y=859900
X3051 4474 2 1 899 BUF1 $T=790500 890520 0 0 $X=790500 $Y=890140
X3052 4545 2 1 4487 BUF1 $T=804760 850200 1 180 $X=802280 $Y=849820
X3053 927 2 1 4381 BUF1 $T=812820 840120 0 180 $X=810340 $Y=834700
X3054 4400 2 1 4666 BUF1 $T=812200 819960 0 0 $X=812200 $Y=819580
X3055 4357 2 1 4676 BUF1 $T=812200 850200 1 0 $X=812200 $Y=844780
X3056 4379 2 1 4700 BUF1 $T=814060 759480 1 0 $X=814060 $Y=754060
X3057 4243 2 1 4710 BUF1 $T=818400 860280 1 0 $X=818400 $Y=854860
X3058 4427 2 1 4720 BUF1 $T=819640 819960 0 0 $X=819640 $Y=819580
X3059 4650 2 1 4739 BUF1 $T=820880 799800 1 0 $X=820880 $Y=794380
X3060 4399 2 1 4721 BUF1 $T=822740 769560 1 0 $X=822740 $Y=764140
X3061 4427 2 1 4736 BUF1 $T=823980 850200 1 0 $X=823980 $Y=844780
X3062 959 2 1 4740 BUF1 $T=837620 739320 0 180 $X=835140 $Y=733900
X3063 4396 2 1 4800 BUF1 $T=835140 759480 1 0 $X=835140 $Y=754060
X3064 4628 2 1 4802 BUF1 $T=835140 799800 1 0 $X=835140 $Y=794380
X3065 4800 2 1 966 BUF1 $T=838860 850200 1 0 $X=838860 $Y=844780
X3066 4824 2 1 967 BUF1 $T=843200 880440 0 180 $X=840720 $Y=875020
X3067 4676 2 1 4819 BUF1 $T=848160 819960 1 180 $X=845680 $Y=819580
X3068 4394 2 1 4863 BUF1 $T=851260 799800 0 0 $X=851260 $Y=799420
X3069 4791 2 1 4912 BUF1 $T=854360 840120 0 0 $X=854360 $Y=839740
X3070 4590 2 1 978 BUF1 $T=856220 880440 0 0 $X=856220 $Y=880060
X3071 987 2 1 4899 BUF1 $T=868000 729240 0 180 $X=865520 $Y=723820
X3072 924 2 1 4953 BUF1 $T=865520 759480 1 0 $X=865520 $Y=754060
X3073 4739 2 1 4968 BUF1 $T=867380 799800 0 0 $X=867380 $Y=799420
X3074 4800 2 1 4918 BUF1 $T=874200 749400 0 0 $X=874200 $Y=749020
X3075 3910 2 1 5010 BUF1 $T=876060 779640 1 0 $X=876060 $Y=774220
X3076 992 2 1 4970 BUF1 $T=884120 870360 0 0 $X=884120 $Y=869980
X3077 4863 2 1 1029 BUF1 $T=899000 809880 0 0 $X=899000 $Y=809500
X3078 4710 2 1 1031 BUF1 $T=901480 880440 1 0 $X=901480 $Y=875020
X3079 5010 2 1 5183 BUF1 $T=903960 809880 0 0 $X=903960 $Y=809500
X3080 5010 2 1 5179 BUF1 $T=905820 759480 0 0 $X=905820 $Y=759100
X3081 1018 2 1 5185 BUF1 $T=906440 809880 1 0 $X=906440 $Y=804460
X3082 992 2 1 1041 BUF1 $T=912020 900600 1 0 $X=912020 $Y=895180
X3083 1038 2 1 5221 BUF1 $T=912640 769560 0 0 $X=912640 $Y=769180
X3084 1020 2 1 5234 BUF1 $T=916980 890520 1 0 $X=916980 $Y=885100
X3085 5221 2 1 1048 BUF1 $T=928760 799800 1 0 $X=928760 $Y=794380
X3086 5257 2 1 5295 BUF1 $T=941160 769560 0 180 $X=938680 $Y=764140
X3087 5356 2 1 1063 BUF1 $T=938680 860280 0 0 $X=938680 $Y=859900
X3088 5257 2 1 5319 BUF1 $T=949840 779640 0 0 $X=949840 $Y=779260
X3089 1025 2 1 1080 BUF1 $T=954180 729240 1 0 $X=954180 $Y=723820
X3090 4361 2 1 5435 BUF1 $T=956040 789720 0 0 $X=956040 $Y=789340
X3091 5307 2 1 1082 BUF1 $T=961620 830040 1 0 $X=961620 $Y=824620
X3092 5528 2 1 5287 BUF1 $T=969060 739320 1 180 $X=966580 $Y=738940
X3093 5385 2 1 5528 BUF1 $T=966580 749400 1 0 $X=966580 $Y=743980
X3094 5557 2 1 1105 BUF1 $T=978980 890520 1 0 $X=978980 $Y=885100
X3095 5687 2 1 5675 BUF1 $T=999440 809880 1 0 $X=999440 $Y=804460
X3096 5704 2 1 5716 BUF1 $T=1004400 739320 0 0 $X=1004400 $Y=738940
X3097 1138 2 1 1115 BUF1 $T=1010600 900600 0 180 $X=1008120 $Y=895180
X3098 1138 2 1 5755 BUF1 $T=1010600 900600 1 0 $X=1010600 $Y=895180
X3099 5663 2 1 1148 BUF1 $T=1014940 779640 0 0 $X=1014940 $Y=779260
X3100 5704 2 1 5749 BUF1 $T=1014940 880440 1 0 $X=1014940 $Y=875020
X3101 5435 2 1 5817 BUF1 $T=1016800 809880 0 0 $X=1016800 $Y=809500
X3102 5749 2 1 1129 BUF1 $T=1019900 890520 1 180 $X=1017420 $Y=890140
X3103 1142 2 1 1153 BUF1 $T=1018040 729240 1 0 $X=1018040 $Y=723820
X3104 5755 2 1 1134 BUF1 $T=1018040 749400 1 0 $X=1018040 $Y=743980
X3105 5689 2 1 1133 BUF1 $T=1020520 880440 1 180 $X=1018040 $Y=880060
X3106 5435 2 1 1147 BUF1 $T=1019280 759480 1 0 $X=1019280 $Y=754060
X3107 5689 2 1 5778 BUF1 $T=1020520 749400 1 0 $X=1020520 $Y=743980
X3108 5649 2 1 5839 BUF1 $T=1021760 809880 1 0 $X=1021760 $Y=804460
X3109 5675 2 1 5855 BUF1 $T=1027960 809880 1 0 $X=1027960 $Y=804460
X3110 5890 2 1 5887 BUF1 $T=1033540 809880 0 0 $X=1033540 $Y=809500
X3111 5935 2 1 1170 BUF1 $T=1039120 739320 1 180 $X=1036640 $Y=738940
X3112 5681 2 1 5924 BUF1 $T=1040360 769560 1 0 $X=1040360 $Y=764140
X3113 5779 2 1 5970 BUF1 $T=1042840 769560 1 0 $X=1042840 $Y=764140
X3114 4976 2 1 1187 BUF1 $T=1045320 819960 0 0 $X=1045320 $Y=819580
X3115 1098 2 1 1192 BUF1 $T=1057720 739320 1 0 $X=1057720 $Y=733900
X3116 1193 2 1 6069 BUF1 $T=1061440 779640 0 0 $X=1061440 $Y=779260
X3117 6018 2 1 6081 BUF1 $T=1064540 809880 0 0 $X=1064540 $Y=809500
X3118 6065 2 1 6047 BUF1 $T=1067020 850200 0 0 $X=1067020 $Y=849820
X3119 1080 2 1 6098 BUF1 $T=1067640 749400 1 0 $X=1067640 $Y=743980
X3120 5855 2 1 6100 BUF1 $T=1068260 819960 1 0 $X=1068260 $Y=814540
X3121 5581 2 1 6122 BUF1 $T=1071360 789720 0 0 $X=1071360 $Y=789340
X3122 1071 2 1 1209 BUF1 $T=1073220 729240 0 0 $X=1073220 $Y=728860
X3123 5840 2 1 1213 BUF1 $T=1076320 890520 0 0 $X=1076320 $Y=890140
X3124 5941 2 1 6147 BUF1 $T=1077560 850200 0 0 $X=1077560 $Y=849820
X3125 5855 2 1 6136 BUF1 $T=1079420 809880 1 0 $X=1079420 $Y=804460
X3126 6150 2 1 6148 BUF1 $T=1080040 850200 0 0 $X=1080040 $Y=849820
X3127 5704 2 1 6162 BUF1 $T=1080660 880440 1 0 $X=1080660 $Y=875020
X3128 1148 2 1 6194 BUF1 $T=1085620 779640 1 0 $X=1085620 $Y=774220
X3129 5581 2 1 6150 BUF1 $T=1089960 830040 1 180 $X=1087480 $Y=829660
X3130 5970 2 1 6248 BUF1 $T=1094920 749400 0 0 $X=1094920 $Y=749020
X3131 6226 2 1 1230 BUF1 $T=1106080 840120 1 180 $X=1103600 $Y=839740
X3132 1213 2 1 6109 BUF1 $T=1105460 890520 1 0 $X=1105460 $Y=885100
X3133 1209 2 1 6293 BUF1 $T=1109800 729240 1 180 $X=1107320 $Y=728860
X3134 6273 2 1 1251 BUF1 $T=1109800 840120 0 0 $X=1109800 $Y=839740
X3135 6293 2 1 6273 BUF1 $T=1114140 789720 1 180 $X=1111660 $Y=789340
X3136 1238 2 1 6065 BUF1 $T=1115380 769560 0 0 $X=1115380 $Y=769180
X3137 6081 2 1 1243 BUF1 $T=1127160 880440 1 180 $X=1124680 $Y=880060
X3138 1520 1 2 1522 BUF1CK $T=254200 840120 0 0 $X=254200 $Y=839740
X3139 1549 1 2 1556 BUF1CK $T=257300 830040 1 0 $X=257300 $Y=824620
X3140 1685 1 2 1692 BUF1CK $T=282720 809880 0 0 $X=282720 $Y=809500
X3141 1704 1 2 1650 BUF1CK $T=287060 789720 1 180 $X=284580 $Y=789340
X3142 1568 1 2 1709 BUF1CK $T=285200 840120 0 0 $X=285200 $Y=839740
X3143 1752 1 2 1765 BUF1CK $T=293260 840120 0 0 $X=293260 $Y=839740
X3144 107 1 2 1764 BUF1CK $T=293880 830040 1 0 $X=293880 $Y=824620
X3145 1772 1 2 1769 BUF1CK $T=296360 830040 1 0 $X=296360 $Y=824620
X3146 1851 1 2 1854 BUF1CK $T=310000 819960 0 0 $X=310000 $Y=819580
X3147 1908 1 2 1915 BUF1CK $T=323020 860280 1 0 $X=323020 $Y=854860
X3148 1911 1 2 1920 BUF1CK $T=323640 840120 1 0 $X=323640 $Y=834700
X3149 136 1 2 1936 BUF1CK $T=326120 860280 0 0 $X=326120 $Y=859900
X3150 2065 1 2 2170 BUF1CK $T=362700 830040 0 0 $X=362700 $Y=829660
X3151 2244 1 2 2248 BUF1CK $T=373240 830040 1 0 $X=373240 $Y=824620
X3152 2236 1 2 2245 BUF1CK $T=376340 840120 0 0 $X=376340 $Y=839740
X3153 1912 1 2 2328 BUF1CK $T=385640 840120 0 0 $X=385640 $Y=839740
X3154 2300 1 2 2528 BUF1CK $T=414780 880440 1 0 $X=414780 $Y=875020
X3155 236 1 2 2521 BUF1CK $T=415400 860280 1 0 $X=415400 $Y=854860
X3156 2641 1 2 2655 BUF1CK $T=440820 779640 1 0 $X=440820 $Y=774220
X3157 276 1 2 2633 BUF1CK $T=440820 860280 0 0 $X=440820 $Y=859900
X3158 2895 1 2 396 BUF1CK $T=491660 880440 0 0 $X=491660 $Y=880060
X3159 3148 1 2 3155 BUF1CK $T=533200 779640 0 0 $X=533200 $Y=779260
X3160 3209 1 2 3214 BUF1CK $T=546840 870360 1 0 $X=546840 $Y=864940
X3161 3262 1 2 3045 BUF1CK $T=559240 779640 0 180 $X=556760 $Y=774220
X3162 481 1 2 3511 BUF1CK $T=598300 900600 1 0 $X=598300 $Y=895180
X3163 2949 1 2 4048 BUF1CK $T=703700 850200 1 0 $X=703700 $Y=844780
X3164 4197 1 2 4235 BUF1CK $T=741520 850200 1 0 $X=741520 $Y=844780
X3165 832 1 2 4328 BUF1CK $T=758880 729240 0 0 $X=758880 $Y=728860
X3166 4337 1 2 4344 BUF1CK $T=759500 890520 1 0 $X=759500 $Y=885100
X3167 4271 1 2 4299 BUF1CK $T=761980 759480 0 0 $X=761980 $Y=759100
X3168 4376 1 2 4519 BUF1CK $T=790500 819960 0 0 $X=790500 $Y=819580
X3169 4636 1 2 4624 BUF1CK $T=807860 789720 1 0 $X=807860 $Y=784300
X3170 932 1 2 4545 BUF1CK $T=815920 890520 0 180 $X=813440 $Y=885100
X3171 4692 1 2 4703 BUF1CK $T=817780 850200 0 0 $X=817780 $Y=849820
X3172 4778 1 2 4776 BUF1CK $T=832660 739320 1 0 $X=832660 $Y=733900
X3173 4857 1 2 4889 BUF1CK $T=855600 860280 1 0 $X=855600 $Y=854860
X3174 4928 1 2 4933 BUF1CK $T=859940 799800 1 0 $X=859940 $Y=794380
X3175 4945 1 2 4946 BUF1CK $T=876680 890520 1 0 $X=876680 $Y=885100
X3176 4914 1 2 4846 BUF1CK $T=879780 890520 0 0 $X=879780 $Y=890140
X3177 4952 1 2 4972 BUF1CK $T=882880 739320 0 0 $X=882880 $Y=738940
X3178 4930 1 2 4835 BUF1CK $T=889080 890520 0 0 $X=889080 $Y=890140
X3179 5138 1 2 5146 BUF1CK $T=898380 739320 0 0 $X=898380 $Y=738940
X3180 5150 1 2 5139 BUF1CK $T=903340 819960 0 0 $X=903340 $Y=819580
X3181 5169 1 2 5187 BUF1CK $T=910780 880440 0 0 $X=910780 $Y=880060
X3182 5274 1 2 5259 BUF1CK $T=926900 769560 1 0 $X=926900 $Y=764140
X3183 5381 1 2 5388 BUF1CK $T=942400 840120 1 0 $X=942400 $Y=834700
X3184 5396 1 2 5407 BUF1CK $T=945500 799800 1 0 $X=945500 $Y=794380
X3185 5459 1 2 5463 BUF1CK $T=954800 830040 0 0 $X=954800 $Y=829660
X3186 5367 1 2 5399 BUF1CK $T=959140 870360 1 0 $X=959140 $Y=864940
X3187 5472 1 2 5503 BUF1CK $T=961000 840120 0 0 $X=961000 $Y=839740
X3188 5513 1 2 5522 BUF1CK $T=964720 830040 1 0 $X=964720 $Y=824620
X3189 5482 1 2 5510 BUF1CK $T=967820 850200 1 0 $X=967820 $Y=844780
X3190 5462 1 2 5439 BUF1CK $T=968440 779640 1 0 $X=968440 $Y=774220
X3191 5560 1 2 5549 BUF1CK $T=972160 749400 0 0 $X=972160 $Y=749020
X3192 5587 1 2 5595 BUF1CK $T=976500 759480 0 0 $X=976500 $Y=759100
X3193 5183 1 2 5581 BUF1CK $T=980840 819960 0 0 $X=980840 $Y=819580
X3194 5637 1 2 5591 BUF1CK $T=984560 850200 0 0 $X=984560 $Y=849820
X3195 5661 1 2 5670 BUF1CK $T=996340 799800 1 0 $X=996340 $Y=794380
X3196 5680 1 2 5688 BUF1CK $T=996960 900600 1 0 $X=996960 $Y=895180
X3197 5648 1 2 5683 BUF1CK $T=998200 819960 0 0 $X=998200 $Y=819580
X3198 5694 1 2 5702 BUF1CK $T=998820 830040 0 0 $X=998820 $Y=829660
X3199 5763 1 2 5771 BUF1CK $T=1007500 830040 0 0 $X=1007500 $Y=829660
X3200 5734 1 2 5695 BUF1CK $T=1008740 850200 0 0 $X=1008740 $Y=849820
X3201 5750 1 2 5759 BUF1CK $T=1009360 769560 0 0 $X=1009360 $Y=769180
X3202 5836 1 2 5834 BUF1CK $T=1022380 809880 0 0 $X=1022380 $Y=809500
X3203 5865 1 2 5871 BUF1CK $T=1026720 799800 0 0 $X=1026720 $Y=799420
X3204 5820 1 2 5804 BUF1CK $T=1029200 749400 1 0 $X=1029200 $Y=743980
X3205 1144 1 2 5890 BUF1CK $T=1029820 860280 1 0 $X=1029820 $Y=854860
X3206 5928 1 2 5937 BUF1CK $T=1036020 819960 0 0 $X=1036020 $Y=819580
X3207 5966 1 2 5962 BUF1CK $T=1043460 809880 1 0 $X=1043460 $Y=804460
X3208 5968 1 2 5969 BUF1CK $T=1044080 729240 0 0 $X=1044080 $Y=728860
X3209 1189 1 2 1190 BUF1CK $T=1049660 890520 0 0 $X=1049660 $Y=890140
X3210 5930 1 2 5903 BUF1CK $T=1057100 890520 1 0 $X=1057100 $Y=885100
X3211 6039 1 2 6030 BUF1CK $T=1059580 850200 0 0 $X=1059580 $Y=849820
X3212 5993 1 2 5950 BUF1CK $T=1072600 870360 1 0 $X=1072600 $Y=864940
X3213 6139 1 2 6121 BUF1CK $T=1078180 759480 1 0 $X=1078180 $Y=754060
X3214 5963 1 2 5917 BUF1CK $T=1078180 860280 0 0 $X=1078180 $Y=859900
X3215 6095 1 2 6118 BUF1CK $T=1081280 749400 0 0 $X=1081280 $Y=749020
X3216 6280 1 2 6247 BUF1CK $T=1107940 880440 0 0 $X=1107940 $Y=880060
X3217 6341 1 2 6330 BUF1CK $T=1112900 870360 0 0 $X=1112900 $Y=869980
X3218 6316 1 2 6367 BUF1CK $T=1114140 890520 0 0 $X=1114140 $Y=890140
X3219 6298 1 2 6295 BUF1CK $T=1114760 819960 0 0 $X=1114760 $Y=819580
X3220 6352 1 2 6370 BUF1CK $T=1125920 840120 0 0 $X=1125920 $Y=839740
X3221 171 1408 1 2 INV2 $T=331700 779640 1 180 $X=329840 $Y=779260
X3222 177 1418 1 2 INV2 $T=332940 789720 1 180 $X=331080 $Y=789340
X3223 174 1955 1 2 INV2 $T=331700 809880 1 0 $X=331700 $Y=804460
X3224 1981 1987 1 2 INV2 $T=333560 789720 0 0 $X=333560 $Y=789340
X3225 2149 2160 1 2 INV2 $T=359600 799800 1 0 $X=359600 $Y=794380
X3226 218 1421 1 2 INV2 $T=361460 749400 0 0 $X=361460 $Y=749020
X3227 2186 2199 1 2 INV2 $T=365800 799800 1 0 $X=365800 $Y=794380
X3228 2214 2234 1 2 INV2 $T=371380 799800 1 0 $X=371380 $Y=794380
X3229 237 1547 1 2 INV2 $T=374480 779640 1 180 $X=372620 $Y=779260
X3230 2260 1704 1 2 INV2 $T=375100 789720 0 180 $X=373240 $Y=784300
X3231 2293 2301 1 2 INV2 $T=381920 789720 1 0 $X=381920 $Y=784300
X3232 253 1500 1 2 INV2 $T=383780 789720 1 0 $X=383780 $Y=784300
X3233 2098 2580 1 2 INV2 $T=426560 789720 0 0 $X=426560 $Y=789340
X3234 2794 2849 1 2 INV2 $T=478640 769560 1 0 $X=478640 $Y=764140
X3235 2655 401 1 2 INV2 $T=492280 749400 1 0 $X=492280 $Y=743980
X3236 2784 2949 1 2 INV2 $T=500340 880440 1 0 $X=500340 $Y=875020
X3237 2580 3248 1 2 INV2 $T=553660 830040 0 0 $X=553660 $Y=829660
X3238 3304 488 1 2 INV2 $T=565440 809880 1 0 $X=565440 $Y=804460
X3239 3448 1690 1 2 INV2 $T=592720 809880 0 180 $X=590860 $Y=804460
X3240 3248 3691 1 2 INV2 $T=642940 830040 1 0 $X=642940 $Y=824620
X3241 3691 3757 1 2 INV2 $T=655340 870360 1 0 $X=655340 $Y=864940
X3242 3352 3859 1 2 INV2 $T=672080 850200 0 0 $X=672080 $Y=849820
X3243 3757 3877 1 2 INV2 $T=675800 840120 0 0 $X=675800 $Y=839740
X3244 4226 420 1 2 INV2 $T=737800 779640 0 0 $X=737800 $Y=779260
X3245 2949 4266 1 2 INV2 $T=745860 850200 1 0 $X=745860 $Y=844780
X3246 4292 686 1 2 INV2 $T=752060 739320 0 180 $X=750200 $Y=733900
X3247 4295 435 1 2 INV2 $T=752060 799800 0 180 $X=750200 $Y=794380
X3248 4318 4309 1 2 INV2 $T=753920 739320 0 0 $X=753920 $Y=738940
X3249 4324 546 1 2 INV2 $T=757640 749400 0 180 $X=755780 $Y=743980
X3250 4222 4276 1 2 INV2 $T=757640 759480 0 0 $X=757640 $Y=759100
X3251 4324 4345 1 2 INV2 $T=759500 749400 0 0 $X=759500 $Y=749020
X3252 812 4334 1 2 INV2 $T=759500 759480 1 0 $X=759500 $Y=754060
X3253 3877 848 1 2 INV2 $T=761980 840120 1 0 $X=761980 $Y=834700
X3254 4284 4271 1 2 INV2 $T=763220 769560 1 0 $X=763220 $Y=764140
X3255 816 4323 1 2 INV2 $T=763840 739320 0 0 $X=763840 $Y=738940
X3256 848 4349 1 2 INV2 $T=764460 840120 1 0 $X=764460 $Y=834700
X3257 4380 839 1 2 INV2 $T=768180 759480 1 0 $X=768180 $Y=754060
X3258 4372 806 1 2 INV2 $T=768180 779640 1 0 $X=768180 $Y=774220
X3259 4348 862 1 2 INV2 $T=771900 769560 1 0 $X=771900 $Y=764140
X3260 4370 888 1 2 INV2 $T=784920 870360 1 0 $X=784920 $Y=864940
X3261 4454 4338 1 2 INV2 $T=786160 809880 1 0 $X=786160 $Y=804460
X3262 4499 4474 1 2 INV2 $T=787400 840120 1 0 $X=787400 $Y=834700
X3263 4578 4485 1 2 INV2 $T=801660 789720 1 180 $X=799800 $Y=789340
X3264 5678 1152 1 2 INV2 $T=1016800 769560 0 0 $X=1016800 $Y=769180
X3265 1152 5779 1 2 INV2 $T=1020520 769560 0 0 $X=1020520 $Y=769180
X3266 6023 6099 1 2 INV2 $T=1068880 809880 1 0 $X=1068880 $Y=804460
X3267 1690 1532 1 2 BUF2 $T=283340 789720 1 180 $X=280240 $Y=789340
X3268 1861 1979 1 2 BUF2 $T=331080 819960 0 0 $X=331080 $Y=819580
X3269 4188 3491 1 2 BUF2 $T=732840 779640 1 180 $X=729740 $Y=779260
X3270 4362 4376 1 2 BUF2 $T=765080 819960 1 0 $X=765080 $Y=814540
X3271 856 3480 1 2 BUF2 $T=769420 779640 1 180 $X=766320 $Y=779260
X3272 4355 865 1 2 BUF2 $T=771900 779640 1 0 $X=771900 $Y=774220
X3273 4517 922 1 2 BUF2 $T=803520 729240 1 0 $X=803520 $Y=723820
X3274 4668 4638 1 2 BUF2 $T=814680 749400 1 0 $X=814680 $Y=743980
X3275 5140 5138 1 2 BUF2 $T=919460 739320 1 0 $X=919460 $Y=733900
X3276 1084 5559 1 2 BUF2 $T=969060 739320 0 0 $X=969060 $Y=738940
X3277 1092 1096 1 2 BUF2 $T=969060 749400 1 0 $X=969060 $Y=743980
X3278 830 5572 1 2 BUF2 $T=971540 769560 1 0 $X=971540 $Y=764140
X3279 5509 5611 1 2 BUF2 $T=978980 819960 1 0 $X=978980 $Y=814540
X3280 806 5644 1 2 BUF2 $T=986420 769560 0 0 $X=986420 $Y=769180
X3281 5606 5560 1 2 BUF2 $T=995720 729240 1 0 $X=995720 $Y=723820
X3282 5936 5991 1 2 BUF2 $T=1046560 789720 0 0 $X=1046560 $Y=789340
X3283 5991 6002 1 2 BUF2 $T=1053380 789720 0 0 $X=1053380 $Y=789340
X3284 5674 1193 1 2 BUF2 $T=1063920 779640 0 0 $X=1063920 $Y=779260
X3285 6299 6341 1 2 BUF2 $T=1106700 840120 0 0 $X=1106700 $Y=839740
X3286 11 1 5 1335 2 1370 ND3 $T=227540 729240 1 0 $X=227540 $Y=723820
X3287 1455 1 1429 1490 2 1483 ND3 $T=247380 870360 1 0 $X=247380 $Y=864940
X3288 1496 1 42 1499 2 45 ND3 $T=249240 880440 0 0 $X=249240 $Y=880060
X3289 1505 1 45 1510 2 1453 ND3 $T=251100 880440 1 0 $X=251100 $Y=875020
X3290 1546 1 53 1492 2 37 ND3 $T=256680 880440 0 180 $X=254200 $Y=875020
X3291 1521 1 1483 1540 2 1453 ND3 $T=256060 870360 1 0 $X=256060 $Y=864940
X3292 1558 1 1607 1596 2 1562 ND3 $T=269080 890520 0 180 $X=266600 $Y=885100
X3293 1512 1 1624 1654 2 1564 ND3 $T=275280 860280 1 0 $X=275280 $Y=854860
X3294 1825 1 1849 1762 2 1796 ND3 $T=309380 890520 0 0 $X=309380 $Y=890140
X3295 125 1 127 1662 2 1856 ND3 $T=310000 870360 1 0 $X=310000 $Y=864940
X3296 1966 1 175 1959 2 1882 ND3 $T=332940 890520 1 180 $X=330460 $Y=890140
X3297 1954 1 1893 1968 2 35 ND3 $T=334800 880440 0 180 $X=332320 $Y=875020
X3298 2166 1 2161 2117 2 2156 ND3 $T=361460 880440 0 180 $X=358980 $Y=875020
X3299 2471 1 2403 2441 2 1796 ND3 $T=408580 880440 1 0 $X=408580 $Y=875020
X3300 2694 1 2688 2682 2 2677 ND3 $T=449500 779640 1 180 $X=447020 $Y=779260
X3301 2701 1 2693 2722 2 2683 ND3 $T=450120 789720 1 0 $X=450120 $Y=784300
X3302 2736 1 2743 2770 2 2733 ND3 $T=461280 799800 1 0 $X=461280 $Y=794380
X3303 2761 1 2754 2769 2 2732 ND3 $T=465000 890520 0 180 $X=462520 $Y=885100
X3304 2774 1 2771 2781 2 2750 ND3 $T=465620 880440 0 180 $X=463140 $Y=875020
X3305 2787 1 2765 2795 2 2783 ND3 $T=467480 789720 1 0 $X=467480 $Y=784300
X3306 2799 1 2805 2814 2 2780 ND3 $T=471200 779640 0 180 $X=468720 $Y=774220
X3307 383 1 2853 385 2 386 ND3 $T=479260 900600 1 0 $X=479260 $Y=895180
X3308 2856 1 2855 2860 2 2858 ND3 $T=480500 789720 1 0 $X=480500 $Y=784300
X3309 2905 1 2903 2914 2 2910 ND3 $T=490420 789720 0 0 $X=490420 $Y=789340
X3310 2918 1 2919 2945 2 2915 ND3 $T=494140 789720 0 0 $X=494140 $Y=789340
X3311 2967 1 2896 2971 2 414 ND3 $T=502200 880440 1 0 $X=502200 $Y=875020
X3312 2983 1 2974 2978 2 2969 ND3 $T=505300 789720 1 180 $X=502820 $Y=789340
X3313 2976 1 2894 2985 2 419 ND3 $T=504060 870360 1 0 $X=504060 $Y=864940
X3314 3006 1 2885 3018 2 3008 ND3 $T=508400 870360 1 0 $X=508400 $Y=864940
X3315 3028 1 2990 3032 2 2980 ND3 $T=512120 880440 0 0 $X=512120 $Y=880060
X3316 3007 1 3050 3058 2 3067 ND3 $T=517700 860280 1 0 $X=517700 $Y=854860
X3317 3072 1 3066 3062 2 3057 ND3 $T=521420 789720 1 180 $X=518940 $Y=789340
X3318 3110 1 3115 3120 2 3111 ND3 $T=527620 880440 1 0 $X=527620 $Y=875020
X3319 3102 1 3113 3108 2 3124 ND3 $T=528240 789720 0 0 $X=528240 $Y=789340
X3320 3133 1 3127 3140 2 439 ND3 $T=531960 870360 1 180 $X=529480 $Y=869980
X3321 3131 1 3136 3138 2 3100 ND3 $T=531340 789720 0 0 $X=531340 $Y=789340
X3322 3416 1 3431 3436 2 3319 ND3 $T=586520 779640 1 0 $X=586520 $Y=774220
X3323 3504 1 3471 3498 2 3197 ND3 $T=601400 890520 0 180 $X=598920 $Y=885100
X3324 3579 1 3583 3611 2 3601 ND3 $T=620620 769560 0 0 $X=620620 $Y=769180
X3325 4018 1 3683 3999 2 718 ND3 $T=700600 769560 1 180 $X=698120 $Y=769180
X3326 4030 1 3643 4016 2 720 ND3 $T=701840 759480 1 180 $X=699360 $Y=759100
X3327 4022 1 3600 4031 2 727 ND3 $T=701220 769560 1 0 $X=701220 $Y=764140
X3328 3229 1 4040 4041 2 4053 ND3 $T=703700 769560 1 0 $X=703700 $Y=764140
X3329 4060 1 3617 4069 2 738 ND3 $T=707420 769560 1 0 $X=707420 $Y=764140
X3330 4078 1 4055 4019 2 733 ND3 $T=709900 840120 1 180 $X=707420 $Y=839740
X3331 4102 1 4085 4044 2 741 ND3 $T=714240 840120 1 180 $X=711760 $Y=839740
X3332 4115 1 4063 4098 2 743 ND3 $T=715480 809880 1 180 $X=713000 $Y=809500
X3333 4164 1 4135 4054 2 764 ND3 $T=727260 809880 1 180 $X=724780 $Y=809500
X3334 4175 1 4150 4042 2 781 ND3 $T=729740 819960 1 0 $X=729740 $Y=814540
X3335 4220 1 4233 4244 2 791 ND3 $T=740280 799800 1 180 $X=737800 $Y=799420
X3336 4314 1 4323 4318 2 4302 ND3 $T=758260 739320 1 180 $X=755780 $Y=738940
X3337 4326 1 4324 603 2 834 ND3 $T=757640 749400 1 0 $X=757640 $Y=743980
X3338 4334 1 4276 837 2 4299 ND3 $T=759500 759480 0 0 $X=759500 $Y=759100
X3339 4323 1 4314 841 2 834 ND3 $T=762600 729240 0 0 $X=762600 $Y=728860
X3340 4222 1 4334 847 2 4271 ND3 $T=764460 759480 1 0 $X=764460 $Y=754060
X3341 4378 1 4389 4174 2 834 ND3 $T=773760 729240 1 180 $X=771280 $Y=728860
X3342 4483 1 4477 4490 2 4473 ND3 $T=786160 809880 0 180 $X=783680 $Y=804460
X3343 4503 1 4500 4509 2 4464 ND3 $T=788020 789720 0 0 $X=788020 $Y=789340
X3344 4520 1 4496 4516 2 4397 ND3 $T=791120 850200 1 180 $X=788640 $Y=849820
X3345 4518 1 4535 4538 2 4419 ND3 $T=794840 789720 1 180 $X=792360 $Y=789340
X3346 4537 1 4524 4547 2 4415 ND3 $T=797320 880440 1 180 $X=794840 $Y=880060
X3347 4577 1 4546 4572 2 4446 ND3 $T=800420 860280 1 180 $X=797940 $Y=859900
X3348 4591 1 916 4602 2 917 ND3 $T=801660 900600 1 0 $X=801660 $Y=895180
X3349 4606 1 4603 4612 2 4429 ND3 $T=806000 799800 0 180 $X=803520 $Y=794380
X3350 4619 1 4593 4627 2 4430 ND3 $T=806620 890520 0 0 $X=806620 $Y=890140
X3351 4732 1 4754 4756 2 4760 ND3 $T=828320 799800 0 0 $X=828320 $Y=799420
X3352 4764 1 4769 4766 2 4783 ND3 $T=831420 759480 1 0 $X=831420 $Y=754060
X3353 4786 1 4775 4613 2 4772 ND3 $T=834520 830040 1 180 $X=832040 $Y=829660
X3354 4879 1 4854 4883 2 4675 ND3 $T=851880 739320 1 180 $X=849400 $Y=738940
X3355 4859 1 4867 4872 2 4874 ND3 $T=849400 759480 1 0 $X=849400 $Y=754060
X3356 4955 1 4957 4947 2 4963 ND3 $T=866760 749400 0 0 $X=866760 $Y=749020
X3357 4929 1 4977 4979 2 4680 ND3 $T=869860 850200 1 0 $X=869860 $Y=844780
X3358 5012 1 5017 5003 2 1001 ND3 $T=877300 870360 0 0 $X=877300 $Y=869980
X3359 5038 1 5041 5032 2 5052 ND3 $T=881640 749400 0 0 $X=881640 $Y=749020
X3360 5064 1 5062 5031 2 1009 ND3 $T=885980 840120 1 180 $X=883500 $Y=839740
X3361 5049 1 5057 5056 2 1012 ND3 $T=883500 860280 0 0 $X=883500 $Y=859900
X3362 5058 1 5073 5077 2 5080 ND3 $T=885980 850200 1 0 $X=885980 $Y=844780
X3363 5078 1 5089 5055 2 1017 ND3 $T=889080 880440 0 0 $X=889080 $Y=880060
X3364 5070 1 5103 5122 2 5111 ND3 $T=891560 749400 0 0 $X=891560 $Y=749020
X3365 5081 1 5145 5175 2 5129 ND3 $T=901480 749400 0 0 $X=901480 $Y=749020
X3366 5088 1 5128 5176 2 5172 ND3 $T=902720 759480 0 0 $X=902720 $Y=759100
X3367 5302 1 5308 5026 2 5318 ND3 $T=931240 749400 0 0 $X=931240 $Y=749020
X3368 5289 1 5311 4521 2 5333 ND3 $T=931240 769560 1 0 $X=931240 $Y=764140
X3369 5303 1 5296 5108 2 5320 ND3 $T=931240 850200 1 0 $X=931240 $Y=844780
X3370 5335 1 1060 4674 2 5359 ND3 $T=937440 880440 0 0 $X=937440 $Y=880060
X3371 5363 1 1062 4689 2 5373 ND3 $T=939920 880440 0 0 $X=939920 $Y=880060
X3372 5370 1 5362 4530 2 5378 ND3 $T=941160 779640 0 0 $X=941160 $Y=779260
X3373 5364 1 5375 5217 2 5382 ND3 $T=941780 759480 1 0 $X=941780 $Y=754060
X3374 5415 1 5395 5067 2 5418 ND3 $T=945500 880440 1 0 $X=945500 $Y=875020
X3375 5397 1 5416 5211 2 5421 ND3 $T=947360 749400 0 0 $X=947360 $Y=749020
X3376 5422 1 5420 4626 2 5406 ND3 $T=949840 779640 1 180 $X=947360 $Y=779260
X3377 5412 1 5369 4595 2 5424 ND3 $T=947360 860280 0 0 $X=947360 $Y=859900
X3378 5417 1 5394 5009 2 5428 ND3 $T=947980 850200 1 0 $X=947980 $Y=844780
X3379 5446 1 5438 5019 2 5458 ND3 $T=952320 850200 0 0 $X=952320 $Y=849820
X3380 5473 1 1083 4686 2 1086 ND3 $T=957900 890520 1 0 $X=957900 $Y=885100
X3381 5484 1 5480 4931 2 5499 ND3 $T=960380 759480 1 0 $X=960380 $Y=754060
X3382 5526 1 5523 5059 2 5511 ND3 $T=967820 850200 0 180 $X=965340 $Y=844780
X3383 5512 1 1090 4618 2 5527 ND3 $T=965340 890520 1 0 $X=965340 $Y=885100
X3384 5488 1 5537 4553 2 5554 ND3 $T=969060 779640 0 0 $X=969060 $Y=779260
X3385 5548 1 5538 4630 2 5558 ND3 $T=970300 880440 1 0 $X=970300 $Y=875020
X3386 5514 1 5563 5114 2 5575 ND3 $T=972160 749400 1 0 $X=972160 $Y=743980
X3387 5515 1 5562 4790 2 5569 ND3 $T=972160 779640 1 0 $X=972160 $Y=774220
X3388 5567 1 5577 4891 2 5594 ND3 $T=975260 739320 0 0 $X=975260 $Y=738940
X3389 5589 1 5565 5033 2 5605 ND3 $T=977120 840120 0 0 $X=977120 $Y=839740
X3390 5601 1 5578 4892 2 5621 ND3 $T=978980 759480 0 0 $X=978980 $Y=759100
X3391 1327 1326 1353 2 1 ND2S $T=222580 840120 1 0 $X=222580 $Y=834700
X3392 1321 1329 1342 2 1 ND2S $T=222580 860280 1 0 $X=222580 $Y=854860
X3393 1340 1353 1367 2 1 ND2S $T=224440 840120 1 0 $X=224440 $Y=834700
X3394 1370 1323 11 2 1 ND2S $T=230020 729240 1 180 $X=228160 $Y=728860
X3395 1348 1342 1307 2 1 ND2S $T=228160 850200 0 0 $X=228160 $Y=849820
X3396 1352 1354 1397 2 1 ND2S $T=231260 860280 1 0 $X=231260 $Y=854860
X3397 1402 1416 1354 2 1 ND2S $T=233740 860280 1 180 $X=231880 $Y=859900
X3398 1370 1423 18 2 1 ND2S $T=236840 729240 1 180 $X=234980 $Y=728860
X3399 19 32 18 2 1 ND2S $T=240560 729240 0 180 $X=238700 $Y=723820
X3400 1432 1451 1431 2 1 ND2S $T=240560 840120 1 180 $X=238700 $Y=839740
X3401 1370 1435 31 2 1 ND2S $T=240560 729240 1 0 $X=240560 $Y=723820
X3402 1472 1489 1451 2 1 ND2S $T=244280 850200 0 180 $X=242420 $Y=844780
X3403 1395 1504 1486 2 1 ND2S $T=247380 819960 0 0 $X=247380 $Y=819580
X3404 1483 1460 1429 2 1 ND2S $T=247380 860280 0 0 $X=247380 $Y=859900
X3405 1492 1479 1499 2 1 ND2S $T=249240 880440 1 180 $X=247380 $Y=880060
X3406 41 39 1483 2 1 ND2S $T=249860 900600 0 180 $X=248000 $Y=895180
X3407 1510 1503 1490 2 1 ND2S $T=252340 870360 0 180 $X=250480 $Y=864940
X3408 1498 1509 1504 2 1 ND2S $T=252960 819960 1 180 $X=251100 $Y=819580
X3409 47 46 1483 2 1 ND2S $T=252960 890520 1 180 $X=251100 $Y=890140
X3410 1449 1511 1522 2 1 ND2S $T=252960 840120 1 0 $X=252960 $Y=834700
X3411 1534 1539 1550 2 1 ND2S $T=256680 809880 0 0 $X=256680 $Y=809500
X3412 1453 1541 1483 2 1 ND2S $T=258540 890520 1 180 $X=256680 $Y=890140
X3413 1525 1550 1347 2 1 ND2S $T=259160 819960 0 180 $X=257300 $Y=814540
X3414 1563 1570 1514 2 1 ND2S $T=261640 809880 1 180 $X=259780 $Y=809500
X3415 1562 1545 1564 2 1 ND2S $T=259780 890520 1 0 $X=259780 $Y=885100
X3416 1485 1571 1518 2 1 ND2S $T=262260 799800 1 180 $X=260400 $Y=799420
X3417 47 65 1564 2 1 ND2S $T=261640 890520 1 0 $X=261640 $Y=885100
X3418 1591 1587 1535 2 1 ND2S $T=269080 870360 0 180 $X=267220 $Y=864940
X3419 1613 1558 47 2 1 ND2S $T=269080 890520 1 0 $X=269080 $Y=885100
X3420 1616 1630 1571 2 1 ND2S $T=272800 809880 0 180 $X=270940 $Y=804460
X3421 1562 1595 1613 2 1 ND2S $T=270940 890520 1 0 $X=270940 $Y=885100
X3422 1636 1640 1570 2 1 ND2S $T=274040 809880 1 0 $X=274040 $Y=804460
X3423 1564 1626 1512 2 1 ND2S $T=274040 860280 0 0 $X=274040 $Y=859900
X3424 1635 1661 72 2 1 ND2S $T=278380 850200 1 180 $X=276520 $Y=849820
X3425 1540 1658 1654 2 1 ND2S $T=279620 860280 0 180 $X=277760 $Y=854860
X3426 1662 1645 1587 2 1 ND2S $T=279620 870360 0 180 $X=277760 $Y=864940
X3427 1612 1696 53 2 1 ND2S $T=283340 850200 1 180 $X=281480 $Y=849820
X3428 1567 1699 1706 2 1 ND2S $T=284580 799800 1 0 $X=284580 $Y=794380
X3429 1719 1707 1699 2 1 ND2S $T=287060 809880 1 180 $X=285200 $Y=809500
X3430 1733 1711 1719 2 1 ND2S $T=290160 799800 0 180 $X=288300 $Y=794380
X3431 1452 1703 1580 2 1 ND2S $T=288300 850200 0 0 $X=288300 $Y=849820
X3432 1712 1742 1678 2 1 ND2S $T=293880 850200 1 180 $X=292020 $Y=849820
X3433 105 1750 1761 2 1 ND2S $T=293880 890520 1 0 $X=293880 $Y=885100
X3434 1750 1676 1762 2 1 ND2S $T=293880 890520 0 0 $X=293880 $Y=890140
X3435 1733 1763 1786 2 1 ND2S $T=295120 809880 1 0 $X=295120 $Y=804460
X3436 1760 1786 1517 2 1 ND2S $T=297600 799800 0 180 $X=295740 $Y=794380
X3437 1794 1800 79 2 1 ND2S $T=300700 850200 0 180 $X=298840 $Y=844780
X3438 1816 1813 1744 2 1 ND2S $T=304420 799800 0 180 $X=302560 $Y=794380
X3439 1802 1780 1813 2 1 ND2S $T=302560 799800 0 0 $X=302560 $Y=799420
X3440 1795 1804 1610 2 1 ND2S $T=302560 809880 0 0 $X=302560 $Y=809500
X3441 1814 1803 109 2 1 ND2S $T=304420 850200 1 180 $X=302560 $Y=849820
X3442 1823 1833 102 2 1 ND2S $T=310000 840120 1 180 $X=308140 $Y=839740
X3443 1612 1852 134 2 1 ND2S $T=310000 850200 0 0 $X=310000 $Y=849820
X3444 1856 1834 127 2 1 ND2S $T=310000 860280 0 0 $X=310000 $Y=859900
X3445 128 123 1849 2 1 ND2S $T=311860 900600 0 180 $X=310000 $Y=895180
X3446 1855 1837 134 2 1 ND2S $T=311860 860280 1 0 $X=311860 $Y=854860
X3447 1635 1863 139 2 1 ND2S $T=313100 850200 0 0 $X=313100 $Y=849820
X3448 1860 1807 1868 2 1 ND2S $T=313100 870360 1 0 $X=313100 $Y=864940
X3449 1452 1880 132 2 1 ND2S $T=316820 850200 0 0 $X=316820 $Y=849820
X3450 1849 1891 149 2 1 ND2S $T=318680 890520 1 180 $X=316820 $Y=890140
X3451 139 1715 153 2 1 ND2S $T=318680 860280 1 0 $X=318680 $Y=854860
X3452 133 1884 1893 2 1 ND2S $T=318680 870360 1 0 $X=318680 $Y=864940
X3453 1886 1870 1882 2 1 ND2S $T=320540 860280 0 0 $X=320540 $Y=859900
X3454 154 1890 132 2 1 ND2S $T=320540 890520 1 0 $X=320540 $Y=885100
X3455 97 1909 1902 2 1 ND2S $T=322400 749400 1 0 $X=322400 $Y=743980
X3456 1613 1896 1512 2 1 ND2S $T=323640 860280 0 0 $X=323640 $Y=859900
X3457 159 1899 1847 2 1 ND2S $T=324260 870360 1 0 $X=324260 $Y=864940
X3458 1564 1927 168 2 1 ND2S $T=326740 870360 1 0 $X=326740 $Y=864940
X3459 1882 1948 168 2 1 ND2S $T=330460 870360 0 180 $X=328600 $Y=864940
X3460 1794 2009 176 2 1 ND2S $T=331080 850200 0 0 $X=331080 $Y=849820
X3461 144 1972 1823 2 1 ND2S $T=332940 860280 0 180 $X=331080 $Y=854860
X3462 1968 1965 1860 2 1 ND2S $T=332940 870360 0 0 $X=332940 $Y=869980
X3463 173 1986 1959 2 1 ND2S $T=336040 900600 0 180 $X=334180 $Y=895180
X3464 1997 2003 1512 2 1 ND2S $T=336660 850200 1 180 $X=334800 $Y=849820
X3465 1882 1989 1512 2 1 ND2S $T=336660 890520 0 180 $X=334800 $Y=885100
X3466 133 1973 2053 2 1 ND2S $T=335420 870360 1 0 $X=335420 $Y=864940
X3467 159 2014 1893 2 1 ND2S $T=337900 880440 0 180 $X=336040 $Y=875020
X3468 1562 2004 1893 2 1 ND2S $T=338520 870360 1 180 $X=336660 $Y=869980
X3469 159 184 1882 2 1 ND2S $T=338520 880440 1 180 $X=336660 $Y=880060
X3470 1996 2008 1712 2 1 ND2S $T=340380 840120 1 180 $X=338520 $Y=839740
X3471 1796 1988 1997 2 1 ND2S $T=338520 860280 1 0 $X=338520 $Y=854860
X3472 1562 2017 1997 2 1 ND2S $T=338520 870360 0 0 $X=338520 $Y=869980
X3473 2073 1991 1984 2 1 ND2S $T=347200 850200 1 0 $X=347200 $Y=844780
X3474 2073 2104 1814 2 1 ND2S $T=352780 850200 1 180 $X=350920 $Y=849820
X3475 1984 2106 209 2 1 ND2S $T=352780 850200 0 0 $X=352780 $Y=849820
X3476 2117 2086 2107 2 1 ND2S $T=352780 880440 1 0 $X=352780 $Y=875020
X3477 2112 2107 2045 2 1 ND2S $T=354640 880440 0 0 $X=354640 $Y=880060
X3478 2122 2126 176 2 1 ND2S $T=358360 850200 0 180 $X=356500 $Y=844780
X3479 144 2123 2151 2 1 ND2S $T=358980 850200 1 0 $X=358980 $Y=844780
X3480 2151 2141 217 2 1 ND2S $T=359600 850200 0 0 $X=359600 $Y=849820
X3481 2156 2136 2161 2 1 ND2S $T=359600 870360 0 0 $X=359600 $Y=869980
X3482 2122 2144 227 2 1 ND2S $T=363940 860280 1 0 $X=363940 $Y=854860
X3483 226 2210 2151 2 1 ND2S $T=368280 819960 1 180 $X=366420 $Y=819580
X3484 153 2183 2211 2 1 ND2S $T=367660 870360 1 0 $X=367660 $Y=864940
X3485 2212 2222 2210 2 1 ND2S $T=369520 809880 1 0 $X=369520 $Y=804460
X3486 2177 2138 2223 2 1 ND2S $T=369520 860280 1 0 $X=369520 $Y=854860
X3487 157 2243 2250 2 1 ND2S $T=375100 819960 0 180 $X=373240 $Y=814540
X3488 2227 2081 2247 2 1 ND2S $T=373240 830040 0 0 $X=373240 $Y=829660
X3489 241 2246 240 2 1 ND2S $T=375720 799800 0 0 $X=375720 $Y=799420
X3490 2257 2278 2227 2 1 ND2S $T=377580 830040 0 0 $X=377580 $Y=829660
X3491 2289 2291 2243 2 1 ND2S $T=381300 819960 0 180 $X=379440 $Y=814540
X3492 2302 2290 2262 2 1 ND2S $T=383160 809880 0 180 $X=381300 $Y=804460
X3493 253 2312 2177 2 1 ND2S $T=384400 799800 0 0 $X=384400 $Y=799420
X3494 2311 2218 2329 2 1 ND2S $T=384400 870360 1 0 $X=384400 $Y=864940
X3495 2342 2351 2312 2 1 ND2S $T=389980 809880 1 180 $X=388120 $Y=809500
X3496 218 2354 1886 2 1 ND2S $T=391220 840120 0 180 $X=389360 $Y=834700
X3497 2311 268 227 2 1 ND2S $T=393700 890520 0 180 $X=391840 $Y=885100
X3498 2382 2369 2354 2 1 ND2S $T=393700 840120 0 0 $X=393700 $Y=839740
X3499 2385 2388 2337 2 1 ND2S $T=394940 809880 0 0 $X=394940 $Y=809500
X3500 274 2406 2074 2 1 ND2S $T=396800 890520 1 180 $X=394940 $Y=890140
X3501 273 2337 2400 2 1 ND2S $T=396800 809880 0 0 $X=396800 $Y=809500
X3502 2330 1947 2403 2 1 ND2S $T=396800 870360 0 0 $X=396800 $Y=869980
X3503 177 2418 2330 2 1 ND2S $T=400520 850200 1 180 $X=398660 $Y=849820
X3504 2396 2419 2418 2 1 ND2S $T=398660 860280 0 0 $X=398660 $Y=859900
X3505 2311 277 2211 2 1 ND2S $T=398660 890520 1 0 $X=398660 $Y=885100
X3506 2447 2416 2433 2 1 ND2S $T=401760 819960 0 0 $X=401760 $Y=819580
X3507 2406 2446 2441 2 1 ND2S $T=402380 880440 1 0 $X=402380 $Y=875020
X3508 171 2436 2397 2 1 ND2S $T=406100 850200 1 0 $X=406100 $Y=844780
X3509 1969 2433 2476 2 1 ND2S $T=407340 830040 0 0 $X=407340 $Y=829660
X3510 2459 2461 2436 2 1 ND2S $T=407340 850200 0 0 $X=407340 $Y=849820
X3511 2397 2477 2420 2 1 ND2S $T=407340 860280 0 0 $X=407340 $Y=859900
X3512 2453 2434 2487 2 1 ND2S $T=409200 840120 1 0 $X=409200 $Y=834700
X3513 237 2487 2506 2 1 ND2S $T=411060 840120 0 0 $X=411060 $Y=839740
X3514 2506 2492 2494 2 1 ND2S $T=412920 850200 1 180 $X=411060 $Y=849820
X3515 1796 2515 2403 2 1 ND2S $T=418500 880440 0 0 $X=418500 $Y=880060
X3516 2699 2694 2643 2 1 ND2S $T=450740 779640 0 180 $X=448880 $Y=774220
X3517 2699 2701 2704 2 1 ND2S $T=449500 779640 0 0 $X=449500 $Y=779260
X3518 2699 2736 2729 2 1 ND2S $T=458800 779640 1 180 $X=456940 $Y=779260
X3519 366 2761 2483 2 1 ND2S $T=464380 880440 1 180 $X=462520 $Y=880060
X3520 366 2774 2778 2 1 ND2S $T=464380 880440 0 0 $X=464380 $Y=880060
X3521 2786 2787 2789 2 1 ND2S $T=466860 779640 0 0 $X=466860 $Y=779260
X3522 2786 2799 2806 2 1 ND2S $T=468720 779640 0 0 $X=468720 $Y=779260
X3523 70 2820 377 2 1 ND2S $T=473060 729240 0 0 $X=473060 $Y=728860
X3524 379 2833 377 2 1 ND2S $T=476780 739320 0 180 $X=474920 $Y=733900
X3525 2786 2856 2818 2 1 ND2S $T=480500 779640 0 0 $X=480500 $Y=779260
X3526 2786 2905 2881 2 1 ND2S $T=491040 789720 1 0 $X=491040 $Y=784300
X3527 2786 2918 2928 2 1 ND2S $T=494760 789720 1 0 $X=494760 $Y=784300
X3528 2923 2967 2847 2 1 ND2S $T=502200 870360 0 0 $X=502200 $Y=869980
X3529 2923 2976 2442 2 1 ND2S $T=504060 870360 0 0 $X=504060 $Y=869980
X3530 2993 2983 2954 2 1 ND2S $T=505300 789720 0 0 $X=505300 $Y=789340
X3531 2923 3006 2897 2 1 ND2S $T=508400 870360 0 180 $X=506540 $Y=864940
X3532 2824 3007 2944 2 1 ND2S $T=510260 860280 1 180 $X=508400 $Y=859900
X3533 2824 3028 3031 2 1 ND2S $T=512120 880440 1 0 $X=512120 $Y=875020
X3534 2993 3072 3056 2 1 ND2S $T=520800 789720 0 180 $X=518940 $Y=784300
X3535 2993 3102 3065 2 1 ND2S $T=523280 789720 0 0 $X=523280 $Y=789340
X3536 2824 3110 3121 2 1 ND2S $T=528240 880440 0 0 $X=528240 $Y=880060
X3537 2824 3133 3078 2 1 ND2S $T=530100 880440 1 0 $X=530100 $Y=875020
X3538 3137 3131 3145 2 1 ND2S $T=531960 789720 1 0 $X=531960 $Y=784300
X3539 3620 3599 3633 2 1 ND2S $T=623100 799800 1 0 $X=623100 $Y=794380
X3540 3619 3630 3631 2 1 ND2S $T=624340 779640 0 0 $X=624340 $Y=779260
X3541 3618 3589 3639 2 1 ND2S $T=626200 779640 1 0 $X=626200 $Y=774220
X3542 3700 3690 3705 2 1 ND2S $T=641080 779640 1 0 $X=641080 $Y=774220
X3543 3893 3878 3770 2 1 ND2S $T=678900 840120 0 180 $X=677040 $Y=834700
X3544 3895 3884 3782 2 1 ND2S $T=680140 850200 1 180 $X=678280 $Y=849820
X3545 3925 3920 3792 2 1 ND2S $T=686340 850200 0 180 $X=684480 $Y=844780
X3546 3922 3957 3813 2 1 ND2S $T=691920 860280 0 180 $X=690060 $Y=854860
X3547 3954 3986 3775 2 1 ND2S $T=695640 819960 1 180 $X=693780 $Y=819580
X3548 4212 4190 4191 2 1 ND2S $T=737180 759480 0 180 $X=735320 $Y=754060
X3549 812 4332 4300 2 1 ND2S $T=760740 779640 0 180 $X=758880 $Y=774220
X3550 4487 4483 4456 2 1 ND2S $T=786160 799800 1 180 $X=784300 $Y=799420
X3551 4497 4506 4492 2 1 ND2S $T=788020 749400 1 180 $X=786160 $Y=749020
X3552 4498 4503 889 2 1 ND2S $T=788020 789720 1 180 $X=786160 $Y=789340
X3553 4532 4525 4440 2 1 ND2S $T=791120 749400 1 180 $X=789260 $Y=749020
X3554 4498 4518 4504 2 1 ND2S $T=791740 799800 0 180 $X=789880 $Y=794380
X3555 4514 4529 4527 2 1 ND2S $T=790500 759480 0 0 $X=790500 $Y=759100
X3556 4545 4537 4536 2 1 ND2S $T=795460 890520 1 180 $X=793600 $Y=890140
X3557 4487 4520 4568 2 1 ND2S $T=799800 850200 0 0 $X=799800 $Y=849820
X3558 913 4591 4452 2 1 ND2S $T=801660 900600 0 180 $X=799800 $Y=895180
X3559 4545 4577 4584 2 1 ND2S $T=801660 870360 1 0 $X=801660 $Y=864940
X3560 4487 4606 4616 2 1 ND2S $T=805380 789720 0 0 $X=805380 $Y=789340
X3561 4545 4619 4601 2 1 ND2S $T=810960 880440 1 180 $X=809100 $Y=880060
X3562 4650 4660 4617 2 1 ND2S $T=814680 799800 1 180 $X=812820 $Y=799420
X3563 4677 4623 4672 2 1 ND2S $T=816540 769560 0 180 $X=814680 $Y=764140
X3564 4628 4659 4714 2 1 ND2S $T=819020 799800 1 0 $X=819020 $Y=794380
X3565 4701 4621 4713 2 1 ND2S $T=819640 840120 1 0 $X=819640 $Y=834700
X3566 4487 4732 4726 2 1 ND2S $T=825840 799800 0 180 $X=823980 $Y=794380
X3567 4743 4684 4748 2 1 ND2S $T=826460 880440 1 0 $X=826460 $Y=875020
X3568 4746 4587 4753 2 1 ND2S $T=827080 870360 1 0 $X=827080 $Y=864940
X3569 4396 4764 4711 2 1 ND2S $T=830180 749400 1 180 $X=828320 $Y=749020
X3570 4752 4667 4758 2 1 ND2S $T=828320 880440 0 0 $X=828320 $Y=880060
X3571 4700 4775 4761 2 1 ND2S $T=833900 830040 0 180 $X=832040 $Y=824620
X3572 4773 4685 4782 2 1 ND2S $T=832040 890520 0 0 $X=832040 $Y=890140
X3573 4700 4769 829 2 1 ND2S $T=833900 749400 0 0 $X=833900 $Y=749020
X3574 4800 4786 4774 2 1 ND2S $T=838860 830040 0 0 $X=838860 $Y=829660
X3575 4871 5024 5023 2 1 ND2S $T=877920 789720 1 0 $X=877920 $Y=784300
X3576 1003 1006 988 2 1 ND2S $T=881640 900600 0 180 $X=879780 $Y=895180
X3577 5030 5025 5039 2 1 ND2S $T=880400 809880 1 0 $X=880400 $Y=804460
X3578 4863 5018 1010 2 1 ND2S $T=881640 799800 1 0 $X=881640 $Y=794380
X3579 1003 5037 4973 2 1 ND2S $T=882260 900600 1 0 $X=882260 $Y=895180
X3580 932 5036 5048 2 1 ND2S $T=887220 890520 0 0 $X=887220 $Y=890140
X3581 4863 5086 5006 2 1 ND2S $T=889080 799800 1 0 $X=889080 $Y=794380
X3582 4871 5106 5060 2 1 ND2S $T=892180 789720 0 180 $X=890320 $Y=784300
X3583 4871 5102 5116 2 1 ND2S $T=892180 789720 0 0 $X=892180 $Y=789340
X3584 4871 5130 5115 2 1 ND2S $T=897760 799800 0 180 $X=895900 $Y=794380
X3585 4863 5131 5120 2 1 ND2S $T=898380 809880 1 180 $X=896520 $Y=809500
X3586 4863 5119 5134 2 1 ND2S $T=899000 799800 1 0 $X=899000 $Y=794380
X3587 4871 5151 5153 2 1 ND2S $T=900860 799800 1 0 $X=900860 $Y=794380
X3588 1029 5159 5165 2 1 ND2S $T=901480 809880 0 0 $X=901480 $Y=809500
X3589 1029 5044 1032 2 1 ND2S $T=901480 890520 0 0 $X=901480 $Y=890140
X3590 5030 5154 5155 2 1 ND2S $T=903340 819960 1 0 $X=903340 $Y=814540
X3591 5030 5091 5193 2 1 ND2S $T=906440 809880 0 0 $X=906440 $Y=809500
X3592 5030 5141 5203 2 1 ND2S $T=908300 809880 0 0 $X=908300 $Y=809500
X3593 5030 5112 5202 2 1 ND2S $T=908920 809880 1 0 $X=908920 $Y=804460
X3594 5706 5752 5732 2 1 ND2S $T=1006260 840120 1 180 $X=1004400 $Y=839740
X3595 5860 5862 5857 2 1 ND2S $T=1027340 850200 0 180 $X=1025480 $Y=844780
X3596 1322 4 1 1322 4 1312 2 MOAI1S $T=223820 880440 1 180 $X=220100 $Y=880060
X3597 1314 1319 1 1314 1319 1332 2 MOAI1S $T=220100 890520 0 0 $X=220100 $Y=890140
X3598 5 1323 1 5 1323 1315 2 MOAI1S $T=224440 749400 0 180 $X=220720 $Y=743980
X3599 1308 1312 1 1308 1312 1337 2 MOAI1S $T=220720 870360 0 0 $X=220720 $Y=869980
X3600 8 1335 1 8 1335 1331 2 MOAI1S $T=226920 729240 0 180 $X=223200 $Y=723820
X3601 9 1341 1 9 1341 1319 2 MOAI1S $T=228160 890520 1 180 $X=224440 $Y=890140
X3602 1368 1369 1 1368 1369 1341 2 MOAI1S $T=231880 900600 0 180 $X=228160 $Y=895180
X3603 1360 1382 1 1360 1382 1386 2 MOAI1S $T=230020 880440 1 0 $X=230020 $Y=875020
X3604 19 1423 1 1398 1376 1343 2 MOAI1S $T=237460 739320 0 180 $X=233740 $Y=733900
X3605 1417 1414 1 1417 1414 1369 2 MOAI1S $T=237460 880440 0 180 $X=233740 $Y=875020
X3606 25 1435 1 28 1443 1444 2 MOAI1S $T=238080 739320 1 0 $X=238080 $Y=733900
X3607 1438 1436 1 1438 1436 1382 2 MOAI1S $T=241800 880440 0 180 $X=238080 $Y=875020
X3608 1457 1456 1 1457 1456 1436 2 MOAI1S $T=245520 880440 0 180 $X=241800 $Y=875020
X3609 1455 1460 1 1455 1460 1469 2 MOAI1S $T=242420 860280 0 0 $X=242420 $Y=859900
X3610 1496 49 1 1496 49 54 2 MOAI1S $T=252960 890520 0 0 $X=252960 $Y=890140
X3611 1437 1537 1 1548 55 1557 2 MOAI1S $T=256060 860280 0 0 $X=256060 $Y=859900
X3612 1533 1544 1 1533 1544 1560 2 MOAI1S $T=256680 880440 0 0 $X=256680 $Y=880060
X3613 1524 1537 1 1548 60 1579 2 MOAI1S $T=257300 830040 0 0 $X=257300 $Y=829660
X3614 1502 1537 1 1548 61 1528 2 MOAI1S $T=258540 850200 0 0 $X=258540 $Y=849820
X3615 1559 1541 1 1559 1541 1314 2 MOAI1S $T=262260 890520 1 180 $X=258540 $Y=890140
X3616 1349 1560 1 1349 1560 1574 2 MOAI1S $T=259160 870360 1 0 $X=259160 $Y=864940
X3617 1338 1537 1 1548 63 1573 2 MOAI1S $T=259780 860280 1 0 $X=259780 $Y=854860
X3618 1551 1537 1 1548 1556 1578 2 MOAI1S $T=262880 830040 1 0 $X=262880 $Y=824620
X3619 1585 66 1 1585 66 1544 2 MOAI1S $T=267220 880440 1 180 $X=263500 $Y=880060
X3620 1333 1537 1 1548 56 1604 2 MOAI1S $T=264120 860280 1 0 $X=264120 $Y=854860
X3621 1600 1596 1 1600 1596 1559 2 MOAI1S $T=268460 890520 1 180 $X=264740 $Y=890140
X3622 1598 1610 1 1615 71 1577 2 MOAI1S $T=267840 819960 1 0 $X=267840 $Y=814540
X3623 1624 1626 1 1624 1626 1632 2 MOAI1S $T=270940 860280 1 0 $X=270940 $Y=854860
X3624 1646 1595 1 1646 1595 1670 2 MOAI1S $T=275900 890520 1 0 $X=275900 $Y=885100
X3625 1674 1610 1 1615 1653 1641 2 MOAI1S $T=280860 819960 1 180 $X=277140 $Y=819580
X3626 1655 82 1 1655 1677 1687 2 MOAI1S $T=279000 729240 0 0 $X=279000 $Y=728860
X3627 1675 1672 1 1675 1672 1456 2 MOAI1S $T=283960 880440 0 180 $X=280240 $Y=875020
X3628 1657 1610 1 1615 1692 1695 2 MOAI1S $T=280860 819960 1 0 $X=280860 $Y=814540
X3629 1658 1693 1 1658 1693 1698 2 MOAI1S $T=282720 860280 1 0 $X=282720 $Y=854860
X3630 1655 93 1 1655 36 96 2 MOAI1S $T=283340 729240 0 0 $X=283340 $Y=728860
X3631 1701 1698 1 1701 1698 1648 2 MOAI1S $T=287060 860280 1 180 $X=283340 $Y=859900
X3632 1723 1721 1 1708 1709 1682 2 MOAI1S $T=288300 840120 0 180 $X=284580 $Y=834700
X3633 1703 1696 1 1703 1696 1718 2 MOAI1S $T=284580 850200 0 0 $X=284580 $Y=849820
X3634 1715 1718 1 1715 1718 1728 2 MOAI1S $T=286440 860280 1 0 $X=286440 $Y=854860
X3635 1745 1721 1 1708 87 1667 2 MOAI1S $T=292640 840120 0 180 $X=288920 $Y=834700
X3636 1661 1728 1 1661 1728 1753 2 MOAI1S $T=290160 860280 1 0 $X=290160 $Y=854860
X3637 1574 1735 1 1574 1735 1748 2 MOAI1S $T=290160 860280 0 0 $X=290160 $Y=859900
X3638 1770 1721 1 1708 91 1747 2 MOAI1S $T=296980 840120 0 180 $X=293260 $Y=834700
X3639 1753 1756 1 1753 1756 1789 2 MOAI1S $T=293880 850200 0 0 $X=293880 $Y=849820
X3640 1758 1748 1 1758 1748 1693 2 MOAI1S $T=297600 860280 1 180 $X=293880 $Y=859900
X3641 1787 1610 1 1615 1769 1757 2 MOAI1S $T=299460 819960 1 180 $X=295740 $Y=819580
X3642 1797 1721 1 1708 1765 1782 2 MOAI1S $T=301320 840120 0 180 $X=297600 $Y=834700
X3643 1791 1789 1 1791 1789 1785 2 MOAI1S $T=301940 860280 0 180 $X=298220 $Y=854860
X3644 1811 1721 1 1708 1793 1799 2 MOAI1S $T=305040 840120 0 180 $X=301320 $Y=834700
X3645 1800 1805 1 1800 1805 1791 2 MOAI1S $T=306280 850200 0 180 $X=302560 $Y=844780
X3646 1807 1803 1 1807 1803 1758 2 MOAI1S $T=306280 860280 1 180 $X=302560 $Y=859900
X3647 1742 1812 1 1742 1812 1831 2 MOAI1S $T=303800 860280 1 0 $X=303800 $Y=854860
X3648 1825 123 1 1825 123 1663 2 MOAI1S $T=309380 900600 0 180 $X=305660 $Y=895180
X3649 1833 1830 1 1833 1830 1805 2 MOAI1S $T=310000 850200 1 180 $X=306280 $Y=849820
X3650 1834 1832 1 1834 1832 1735 2 MOAI1S $T=310000 860280 1 180 $X=306280 $Y=859900
X3651 1837 1831 1 1837 1831 1756 2 MOAI1S $T=311240 860280 0 180 $X=307520 $Y=854860
X3652 1746 1828 1 1843 1777 1876 2 MOAI1S $T=311240 830040 1 0 $X=311240 $Y=824620
X3653 1809 1865 1 141 1872 1877 2 MOAI1S $T=313100 739320 1 0 $X=313100 $Y=733900
X3654 1870 1867 1 1870 1867 1792 2 MOAI1S $T=317440 860280 0 180 $X=313720 $Y=854860
X3655 1884 1883 1 1884 1883 1832 2 MOAI1S $T=320540 860280 1 180 $X=316820 $Y=859900
X3656 1891 1890 1 1891 1890 1812 2 MOAI1S $T=322400 880440 1 180 $X=318680 $Y=880060
X3657 1899 1896 1 1899 1896 1883 2 MOAI1S $T=324260 870360 0 180 $X=320540 $Y=864940
X3658 1943 1844 1 1926 1915 1905 2 MOAI1S $T=329220 850200 0 180 $X=325500 $Y=844780
X3659 1927 1923 1 1927 1923 1867 2 MOAI1S $T=329220 860280 0 180 $X=325500 $Y=854860
X3660 1949 1942 1 1829 1920 1907 2 MOAI1S $T=329840 840120 0 180 $X=326120 $Y=834700
X3661 169 1952 1 1940 1901 1931 2 MOAI1S $T=331080 739320 0 180 $X=327360 $Y=733900
X3662 1958 1844 1 1926 165 1925 2 MOAI1S $T=331080 840120 1 180 $X=327360 $Y=839740
X3663 170 1952 1 1940 1944 1898 2 MOAI1S $T=331700 749400 1 180 $X=327980 $Y=749020
X3664 1933 1942 1 1945 1941 1939 2 MOAI1S $T=331700 799800 0 180 $X=327980 $Y=794380
X3665 1918 1942 1 1945 1919 1932 2 MOAI1S $T=331700 809880 0 180 $X=327980 $Y=804460
X3666 1938 1942 1 1945 1961 1906 2 MOAI1S $T=328600 799800 0 0 $X=328600 $Y=799420
X3667 1863 1947 1 1863 1947 1964 2 MOAI1S $T=328600 860280 0 0 $X=328600 $Y=859900
X3668 1971 1844 1 1829 1773 1956 2 MOAI1S $T=333560 840120 0 180 $X=329840 $Y=834700
X3669 1980 1844 1 1926 1936 1946 2 MOAI1S $T=333560 850200 0 180 $X=329840 $Y=844780
X3670 1973 1964 1 1973 1964 1998 2 MOAI1S $T=332940 860280 0 0 $X=332940 $Y=859900
X3671 1991 1988 1 1991 1988 1923 2 MOAI1S $T=337900 860280 0 180 $X=334180 $Y=854860
X3672 1966 1989 1 1966 1989 2018 2 MOAI1S $T=334180 890520 0 0 $X=334180 $Y=890140
X3673 2030 1942 1 1945 1979 1985 2 MOAI1S $T=340380 819960 1 180 $X=336660 $Y=819580
X3674 2004 1998 1 2004 1998 2023 2 MOAI1S $T=336660 860280 0 0 $X=336660 $Y=859900
X3675 1937 1942 1 1945 2022 2025 2 MOAI1S $T=337280 809880 0 0 $X=337280 $Y=809500
X3676 2003 2008 1 2003 2008 2031 2 MOAI1S $T=337280 850200 1 0 $X=337280 $Y=844780
X3677 2009 2015 1 2009 2015 2037 2 MOAI1S $T=337900 850200 0 0 $X=337900 $Y=849820
X3678 2023 2034 1 2023 2034 2047 2 MOAI1S $T=340380 860280 1 0 $X=340380 $Y=854860
X3679 1967 2038 1 1967 2038 2060 2 MOAI1S $T=341000 870360 0 0 $X=341000 $Y=869980
X3680 1880 2037 1 1880 2037 2059 2 MOAI1S $T=342240 850200 0 0 $X=342240 $Y=849820
X3681 2059 2047 1 2059 2047 2041 2 MOAI1S $T=347820 860280 0 180 $X=344100 $Y=854860
X3682 1852 2072 1 1852 2072 2085 2 MOAI1S $T=346580 850200 0 0 $X=346580 $Y=849820
X3683 2081 2031 1 2081 2031 2072 2 MOAI1S $T=350920 840120 1 180 $X=347200 $Y=839740
X3684 2082 2077 1 2082 2077 2038 2 MOAI1S $T=350920 860280 1 180 $X=347200 $Y=859900
X3685 2090 2085 1 2090 2085 2034 2 MOAI1S $T=352160 860280 0 180 $X=348440 $Y=854860
X3686 2111 2105 1 2111 2105 2077 2 MOAI1S $T=354640 870360 0 180 $X=350920 $Y=864940
X3687 1953 2106 1 1953 2106 2082 2 MOAI1S $T=354640 870360 1 180 $X=350920 $Y=869980
X3688 2119 2104 1 2119 2104 2111 2 MOAI1S $T=355880 860280 0 180 $X=352160 $Y=854860
X3689 2126 2123 1 2126 2123 1830 2 MOAI1S $T=356500 850200 0 180 $X=352780 $Y=844780
X3690 2148 2063 1 2007 151 2069 2 MOAI1S $T=357740 840120 1 180 $X=354020 $Y=839740
X3691 2136 2135 1 2136 2135 2090 2 MOAI1S $T=358360 870360 0 180 $X=354640 $Y=864940
X3692 2141 2138 1 2141 2138 2015 2 MOAI1S $T=358980 850200 1 180 $X=355260 $Y=849820
X3693 2147 2144 1 2147 2144 2119 2 MOAI1S $T=359600 860280 1 180 $X=355880 $Y=859900
X3694 2139 2055 1 2139 2055 2158 2 MOAI1S $T=356500 880440 0 0 $X=356500 $Y=880060
X3695 2165 2063 1 2007 2153 2110 2 MOAI1S $T=361460 840120 1 180 $X=357740 $Y=839740
X3696 214 1972 1 214 1972 2147 2 MOAI1S $T=362080 860280 0 180 $X=358360 $Y=854860
X3697 2093 1828 1 2058 2170 2174 2 MOAI1S $T=358980 830040 0 0 $X=358980 $Y=829660
X3698 2140 224 1 2140 224 2197 2 MOAI1S $T=363320 890520 0 0 $X=363320 $Y=890140
X3699 2183 1948 1 2183 1948 2208 2 MOAI1S $T=364560 860280 0 0 $X=364560 $Y=859900
X3700 2215 1828 1 2058 2189 2185 2 MOAI1S $T=368900 830040 1 180 $X=365180 $Y=829660
X3701 2218 2208 1 2218 2208 2135 2 MOAI1S $T=372620 860280 1 180 $X=368900 $Y=859900
X3702 2252 2246 1 241 240 2217 2 MOAI1S $T=375720 799800 1 180 $X=372000 $Y=799420
X3703 246 2063 1 2007 2245 2240 2 MOAI1S $T=376960 850200 0 180 $X=373240 $Y=844780
X3704 2295 2063 1 2007 247 2229 2 MOAI1S $T=382540 840120 1 180 $X=378820 $Y=839740
X3705 2296 2063 1 2007 203 2195 2 MOAI1S $T=382540 850200 0 180 $X=378820 $Y=844780
X3706 2271 2288 1 2271 2288 2292 2 MOAI1S $T=380060 890520 1 0 $X=380060 $Y=885100
X3707 2158 2292 1 2158 2292 2315 2 MOAI1S $T=380680 880440 0 0 $X=380680 $Y=880060
X3708 2304 2268 1 2304 2268 2320 2 MOAI1S $T=382540 870360 0 0 $X=382540 $Y=869980
X3709 2340 2334 1 2058 255 2253 2 MOAI1S $T=387500 830040 1 180 $X=383780 $Y=829660
X3710 2350 2334 1 2325 172 2314 2 MOAI1S $T=388120 850200 0 180 $X=384400 $Y=844780
X3711 2307 2334 1 2325 2328 2316 2 MOAI1S $T=388740 840120 0 180 $X=385020 $Y=834700
X3712 2320 2315 1 2320 2315 2344 2 MOAI1S $T=385020 880440 0 0 $X=385020 $Y=880060
X3713 2324 2343 1 2325 2248 2327 2 MOAI1S $T=389360 830040 0 180 $X=385640 $Y=824620
X3714 2356 190 1 1843 2319 2332 2 MOAI1S $T=390600 870360 1 180 $X=386880 $Y=869980
X3715 2197 2344 1 2197 2344 266 2 MOAI1S $T=388120 890520 1 0 $X=388120 $Y=885100
X3716 2311 2161 1 2310 252 263 2 MOAI1S $T=393700 880440 1 180 $X=389980 $Y=880060
X3717 2391 190 1 1843 270 2348 2 MOAI1S $T=396180 870360 1 180 $X=392460 $Y=869980
X3718 2378 2343 1 2325 2390 2393 2 MOAI1S $T=393080 830040 0 0 $X=393080 $Y=829660
X3719 2381 2343 1 2325 2235 2395 2 MOAI1S $T=393700 819960 0 0 $X=393700 $Y=819580
X3720 2386 2334 1 2325 249 2402 2 MOAI1S $T=394940 850200 1 0 $X=394940 $Y=844780
X3721 2311 2223 1 249 276 278 2 MOAI1S $T=395560 880440 1 0 $X=395560 $Y=875020
X3722 2492 2477 1 2492 2477 2105 2 MOAI1S $T=413540 860280 1 180 $X=409820 $Y=859900
X3723 2471 2515 1 2471 2515 2529 2 MOAI1S $T=414160 880440 0 0 $X=414160 $Y=880060
X3724 299 2530 1 2522 2521 2496 2 MOAI1S $T=418500 870360 0 180 $X=414780 $Y=864940
X3725 305 2530 1 2522 2219 2512 2 MOAI1S $T=422220 870360 0 180 $X=418500 $Y=864940
X3726 308 2530 1 2522 2528 2555 2 MOAI1S $T=426560 870360 1 180 $X=422840 $Y=869980
X3727 314 2530 1 2546 2095 2562 2 MOAI1S $T=428420 860280 1 180 $X=424700 $Y=859900
X3728 318 2571 1 2546 2134 2572 2 MOAI1S $T=430280 850200 0 180 $X=426560 $Y=844780
X3729 2589 2554 1 1940 2377 2567 2 MOAI1S $T=430900 809880 1 180 $X=427180 $Y=809500
X3730 322 2554 1 1940 2519 2578 2 MOAI1S $T=431520 819960 0 180 $X=427800 $Y=814540
X3731 2599 2554 1 2546 2318 2582 2 MOAI1S $T=432760 840120 0 180 $X=429040 $Y=834700
X3732 324 2571 1 2546 2190 2592 2 MOAI1S $T=434620 850200 0 180 $X=430900 $Y=844780
X3733 327 2571 1 2522 2603 2606 2 MOAI1S $T=437100 870360 0 180 $X=433380 $Y=864940
X3734 334 2571 1 2522 2633 2629 2 MOAI1S $T=441440 870360 0 180 $X=437720 $Y=864940
X3735 2841 2439 1 2670 2857 2752 2 MOAI1S $T=478020 809880 0 0 $X=478020 $Y=809500
X3736 2773 2893 1 2773 2857 2844 2 MOAI1S $T=489180 850200 0 180 $X=485460 $Y=844780
X3737 2717 397 1 2717 399 2912 2 MOAI1S $T=489180 870360 0 0 $X=489180 $Y=869980
X3738 2866 2917 1 2866 2857 2901 2 MOAI1S $T=494760 830040 0 180 $X=491040 $Y=824620
X3739 2845 2913 1 2845 2857 2922 2 MOAI1S $T=491660 830040 0 0 $X=491660 $Y=829660
X3740 2937 2948 1 2937 2857 2900 2 MOAI1S $T=500340 809880 0 180 $X=496620 $Y=804460
X3741 2773 2384 1 2773 399 2955 2 MOAI1S $T=496620 860280 1 0 $X=496620 $Y=854860
X3742 394 2950 1 394 404 2932 2 MOAI1S $T=500340 900600 0 180 $X=496620 $Y=895180
X3743 2956 2959 1 2956 399 2946 2 MOAI1S $T=500340 870360 1 0 $X=500340 $Y=864940
X3744 2876 2972 1 2977 2987 2991 2 MOAI1S $T=502820 779640 0 0 $X=502820 $Y=779260
X3745 2956 2973 1 2956 415 2975 2 MOAI1S $T=507780 860280 1 180 $X=504060 $Y=859900
X3746 2999 3011 1 2956 3003 2995 2 MOAI1S $T=510880 880440 0 180 $X=507160 $Y=875020
X3747 2866 3005 1 2866 3003 3020 2 MOAI1S $T=507780 830040 0 0 $X=507780 $Y=829660
X3748 2965 3038 1 2965 3003 3017 2 MOAI1S $T=515840 819960 1 180 $X=512120 $Y=819580
X3749 403 3030 1 403 399 3040 2 MOAI1S $T=512120 900600 1 0 $X=512120 $Y=895180
X3750 3068 2573 1 380 404 3046 2 MOAI1S $T=520800 880440 1 180 $X=517080 $Y=880060
X3751 3093 3104 1 3093 3092 3081 2 MOAI1S $T=527620 819960 1 180 $X=523900 $Y=819580
X3752 2882 2423 1 2882 3092 3083 2 MOAI1S $T=529480 860280 0 180 $X=525760 $Y=854860
X3753 2999 3142 1 2999 446 3150 2 MOAI1S $T=531960 880440 0 0 $X=531960 $Y=880060
X3754 3095 443 1 3095 446 3158 2 MOAI1S $T=531960 890520 0 0 $X=531960 $Y=890140
X3755 3149 3155 1 3149 2987 3143 2 MOAI1S $T=536920 779640 0 180 $X=533200 $Y=774220
X3756 2937 2408 1 2937 3161 3164 2 MOAI1S $T=533200 809880 1 0 $X=533200 $Y=804460
X3757 2999 3130 1 2999 447 3166 2 MOAI1S $T=533200 880440 1 0 $X=533200 $Y=875020
X3758 2977 3156 1 2977 3167 3171 2 MOAI1S $T=534440 789720 1 0 $X=534440 $Y=784300
X3759 2965 3152 1 2965 3092 3175 2 MOAI1S $T=535060 830040 1 0 $X=535060 $Y=824620
X3760 3004 3014 1 3004 3092 3172 2 MOAI1S $T=541260 809880 0 180 $X=537540 $Y=804460
X3761 3068 3178 1 3068 3189 3194 2 MOAI1S $T=538780 860280 1 0 $X=538780 $Y=854860
X3762 3215 3226 1 3215 415 3203 2 MOAI1S $T=551800 819960 1 180 $X=548080 $Y=819580
X3763 466 469 1 466 3189 3195 2 MOAI1S $T=554900 870360 1 180 $X=551180 $Y=869980
X3764 3247 3255 1 3247 3248 3231 2 MOAI1S $T=557380 840120 1 180 $X=553660 $Y=839740
X3765 3061 3258 1 3061 2987 3230 2 MOAI1S $T=558620 769560 1 180 $X=554900 $Y=769180
X3766 3256 3224 1 3061 3263 3261 2 MOAI1S $T=561100 779640 1 180 $X=557380 $Y=779260
X3767 3247 3277 1 3247 3151 3303 2 MOAI1S $T=559240 819960 0 0 $X=559240 $Y=819580
X3768 3271 2520 1 3271 3189 3251 2 MOAI1S $T=562960 870360 0 180 $X=559240 $Y=864940
X3769 3287 3293 1 3215 3151 3308 2 MOAI1S $T=562340 840120 1 0 $X=562340 $Y=834700
X3770 3204 3325 1 3204 2987 3311 2 MOAI1S $T=569780 749400 1 180 $X=566060 $Y=749020
X3771 3332 3344 1 3332 3250 3327 2 MOAI1S $T=571020 799800 1 0 $X=571020 $Y=794380
X3772 3252 3039 1 3252 2987 3367 2 MOAI1S $T=574120 749400 0 0 $X=574120 $Y=749020
X3773 3256 3383 1 3256 507 3365 2 MOAI1S $T=579700 789720 0 180 $X=575980 $Y=784300
X3774 506 509 1 506 507 514 2 MOAI1S $T=576600 729240 0 0 $X=576600 $Y=728860
X3775 3345 510 1 3345 3248 3405 2 MOAI1S $T=576600 819960 0 0 $X=576600 $Y=819580
X3776 511 3337 1 3370 3250 3371 2 MOAI1S $T=581560 880440 0 180 $X=577840 $Y=875020
X3777 3382 513 1 3382 3407 3388 2 MOAI1S $T=578460 739320 0 0 $X=578460 $Y=738940
X3778 3382 3391 1 3382 507 3411 2 MOAI1S $T=578460 749400 1 0 $X=578460 $Y=743980
X3779 3370 2352 1 3370 3189 3421 2 MOAI1S $T=581560 870360 0 0 $X=581560 $Y=869980
X3780 506 521 1 506 529 3425 2 MOAI1S $T=583420 729240 0 0 $X=583420 $Y=728860
X3781 524 527 1 524 529 3435 2 MOAI1S $T=584660 739320 1 0 $X=584660 $Y=733900
X3782 3432 3427 1 3432 3248 3437 2 MOAI1S $T=587140 830040 0 0 $X=587140 $Y=829660
X3783 3413 3439 1 3413 3225 3396 2 MOAI1S $T=591480 769560 0 180 $X=587760 $Y=764140
X3784 3332 2640 1 3332 3393 3444 2 MOAI1S $T=588380 789720 1 0 $X=588380 $Y=784300
X3785 3332 539 1 3332 3463 3451 2 MOAI1S $T=592720 789720 0 0 $X=592720 $Y=789340
X3786 3501 3477 1 3428 3189 3479 2 MOAI1S $T=601400 860280 1 180 $X=597680 $Y=859900
X3787 3485 2608 1 3485 3189 3476 2 MOAI1S $T=601400 870360 0 180 $X=597680 $Y=864940
X3788 3464 3509 1 3464 3520 3524 2 MOAI1S $T=601400 840120 1 0 $X=601400 $Y=834700
X3789 3464 3366 1 3464 3248 3535 2 MOAI1S $T=603880 830040 0 0 $X=603880 $Y=829660
X3790 3485 3530 1 3464 3536 3540 2 MOAI1S $T=604500 860280 1 0 $X=604500 $Y=854860
X3791 3527 555 1 3527 537 3496 2 MOAI1S $T=609460 749400 1 180 $X=605740 $Y=749020
X3792 3546 3543 1 554 3250 3531 2 MOAI1S $T=610080 890520 0 180 $X=606360 $Y=885100
X3793 3501 3542 1 3501 3248 3558 2 MOAI1S $T=608220 830040 0 0 $X=608220 $Y=829660
X3794 3554 564 1 3554 537 3526 2 MOAI1S $T=615040 759480 0 180 $X=611320 $Y=754060
X3795 3428 559 1 3428 3536 3556 2 MOAI1S $T=611320 860280 1 0 $X=611320 $Y=854860
X3796 3527 3567 1 3527 3407 3541 2 MOAI1S $T=616280 739320 1 180 $X=612560 $Y=738940
X3797 563 2581 1 563 3250 3557 2 MOAI1S $T=616280 890520 0 180 $X=612560 $Y=885100
X3798 3563 3570 1 3563 537 3537 2 MOAI1S $T=616900 779640 0 180 $X=613180 $Y=774220
X3799 565 3499 1 565 3407 3505 2 MOAI1S $T=617520 729240 1 180 $X=613800 $Y=728860
X3800 3554 3565 1 3554 3407 3576 2 MOAI1S $T=620620 739320 1 180 $X=616900 $Y=738940
X3801 3528 573 1 3584 537 3538 2 MOAI1S $T=620620 779640 0 180 $X=616900 $Y=774220
X3802 3584 2666 1 3528 3263 3539 2 MOAI1S $T=618140 789720 1 0 $X=618140 $Y=784300
X3803 3501 2621 1 3501 3597 3605 2 MOAI1S $T=618140 840120 1 0 $X=618140 $Y=834700
X3804 3549 3580 1 3549 3263 3550 2 MOAI1S $T=623100 799800 0 180 $X=619380 $Y=794380
X3805 578 580 1 578 3407 588 2 MOAI1S $T=623720 729240 0 0 $X=623720 $Y=728860
X3806 3527 583 1 3606 589 3598 2 MOAI1S $T=624340 739320 0 0 $X=624340 $Y=738940
X3807 3563 3632 1 3563 3263 3645 2 MOAI1S $T=624960 789720 0 0 $X=624960 $Y=789340
X3808 3606 594 1 3606 534 3674 2 MOAI1S $T=629300 739320 0 0 $X=629300 $Y=738940
X3809 597 3640 1 597 589 3681 2 MOAI1S $T=632400 729240 0 0 $X=632400 $Y=728860
X3810 3662 3665 1 3662 3463 3685 2 MOAI1S $T=633020 749400 0 0 $X=633020 $Y=749020
X3811 3678 3642 1 3563 3463 3663 2 MOAI1S $T=636740 779640 0 180 $X=633020 $Y=774220
X3812 3693 617 1 3693 3664 3721 2 MOAI1S $T=639220 819960 1 0 $X=639220 $Y=814540
X3813 3637 3624 1 3697 3686 3613 2 MOAI1S $T=643560 809880 0 180 $X=639840 $Y=804460
X3814 3669 623 1 3655 3664 3672 2 MOAI1S $T=643560 870360 1 180 $X=639840 $Y=869980
X3815 3528 2698 1 3706 3714 3731 2 MOAI1S $T=642940 789720 0 0 $X=642940 $Y=789340
X3816 3549 3719 1 3549 3714 3716 2 MOAI1S $T=646660 799800 1 180 $X=642940 $Y=799420
X3817 3737 3762 1 3737 3536 3717 2 MOAI1S $T=654720 850200 0 180 $X=651000 $Y=844780
X3818 3729 3615 1 3729 3757 3722 2 MOAI1S $T=655340 870360 0 180 $X=651620 $Y=864940
X3819 3737 3807 1 3737 3714 3789 2 MOAI1S $T=662780 840120 0 180 $X=659060 $Y=834700
X3820 3825 662 1 3825 3757 3783 2 MOAI1S $T=668360 870360 0 180 $X=664640 $Y=864940
X3821 3858 3310 1 3858 3597 3840 2 MOAI1S $T=675800 840120 1 180 $X=672080 $Y=839740
X3822 3858 3725 1 3858 3757 3853 2 MOAI1S $T=679520 870360 0 180 $X=675800 $Y=864940
X3823 3956 712 1 3956 3714 3993 2 MOAI1S $T=693160 850200 1 0 $X=693160 $Y=844780
X3824 4127 753 1 4127 4136 4140 2 MOAI1S $T=717340 830040 0 0 $X=717340 $Y=829660
X3825 4159 769 1 4159 3714 4158 2 MOAI1S $T=728500 840120 1 180 $X=724780 $Y=839740
X3826 4159 4142 1 4159 4167 4165 2 MOAI1S $T=725400 860280 1 0 $X=725400 $Y=854860
X3827 4180 4213 1 4180 4167 4177 2 MOAI1S $T=737800 860280 0 180 $X=734080 $Y=854860
X3828 4191 768 1 4201 4229 792 2 MOAI1S $T=735940 749400 1 0 $X=735940 $Y=743980
X3829 4180 4235 1 4180 4243 4245 2 MOAI1S $T=738420 860280 1 0 $X=738420 $Y=854860
X3830 4234 4237 1 4234 4136 4254 2 MOAI1S $T=739040 819960 0 0 $X=739040 $Y=819580
X3831 4176 4238 1 4176 4136 4269 2 MOAI1S $T=739040 830040 1 0 $X=739040 $Y=824620
X3832 4264 4273 1 4264 4243 4283 2 MOAI1S $T=745860 860280 1 0 $X=745860 $Y=854860
X3833 4264 821 1 4264 3859 4296 2 MOAI1S $T=748340 860280 0 0 $X=748340 $Y=859900
X3834 4359 4344 1 838 4338 4287 2 MOAI1S $T=763220 890520 1 180 $X=759500 $Y=890140
X3835 4360 850 1 4360 4136 4297 2 MOAI1S $T=767560 809880 0 180 $X=763840 $Y=804460
X3836 4360 851 1 4360 4361 4298 2 MOAI1S $T=768180 809880 1 180 $X=764460 $Y=809500
X3837 4352 4371 1 4352 4338 4354 2 MOAI1S $T=768180 890520 0 180 $X=764460 $Y=885100
X3838 4374 4363 1 4374 4370 4364 2 MOAI1S $T=770040 860280 1 180 $X=766320 $Y=859900
X3839 838 4398 1 838 848 4340 2 MOAI1S $T=772520 890520 1 180 $X=768800 $Y=890140
X3840 4391 860 1 4391 4361 4321 2 MOAI1S $T=773140 799800 1 180 $X=769420 $Y=799420
X3841 4352 4281 1 4352 4370 4375 2 MOAI1S $T=776240 860280 1 180 $X=772520 $Y=859900
X3842 4391 4436 1 4391 4136 4417 2 MOAI1S $T=777480 809880 0 180 $X=773760 $Y=804460
X3843 4422 4449 1 4422 4434 4426 2 MOAI1S $T=779340 769560 1 180 $X=775620 $Y=769180
X3844 4407 877 1 4407 4437 4405 2 MOAI1S $T=780580 830040 1 180 $X=776860 $Y=829660
X3845 4450 4460 1 4450 4437 4421 2 MOAI1S $T=782440 819960 0 180 $X=778720 $Y=814540
X3846 4455 4457 1 4455 4434 4476 2 MOAI1S $T=779960 759480 1 0 $X=779960 $Y=754060
X3847 4448 4484 1 4448 881 4441 2 MOAI1S $T=786160 789720 1 180 $X=782440 $Y=789340
X3848 4491 893 1 4491 4480 4459 2 MOAI1S $T=788640 860280 1 180 $X=784920 $Y=859900
X3849 4491 4432 1 4491 4338 4413 2 MOAI1S $T=788640 880440 1 180 $X=784920 $Y=880060
X3850 4422 891 1 4422 881 4469 2 MOAI1S $T=786160 759480 0 0 $X=786160 $Y=759100
X3851 4455 895 1 4455 881 4489 2 MOAI1S $T=787400 749400 1 0 $X=787400 $Y=743980
X3852 4448 4507 1 4448 4517 4515 2 MOAI1S $T=788020 789720 1 0 $X=788020 $Y=784300
X3853 4512 901 1 4512 4480 4549 2 MOAI1S $T=792360 870360 1 0 $X=792360 $Y=864940
X3854 4455 4543 1 4455 4517 4562 2 MOAI1S $T=794220 749400 0 0 $X=794220 $Y=749020
X3855 4544 4550 1 4544 906 4569 2 MOAI1S $T=794840 890520 1 0 $X=794840 $Y=885100
X3856 4575 909 1 4422 4517 4558 2 MOAI1S $T=799800 759480 1 180 $X=796080 $Y=759100
X3857 4566 908 1 4566 4517 4557 2 MOAI1S $T=797940 739320 1 0 $X=797940 $Y=733900
X3858 4566 4570 1 4566 4434 4552 2 MOAI1S $T=797940 739320 0 0 $X=797940 $Y=738940
X3859 4580 915 1 4580 4517 4573 2 MOAI1S $T=803520 729240 0 180 $X=799800 $Y=723820
X3860 4560 4528 1 4560 4361 4609 2 MOAI1S $T=801660 830040 0 0 $X=801660 $Y=829660
X3861 4566 4607 1 4566 881 4592 2 MOAI1S $T=806000 739320 1 180 $X=802280 $Y=738940
X3862 4596 4610 1 4596 4480 4635 2 MOAI1S $T=804140 860280 0 0 $X=804140 $Y=859900
X3863 4580 4638 1 4580 4434 4620 2 MOAI1S $T=810340 739320 0 180 $X=806620 $Y=733900
X3864 4608 4624 1 4608 4338 4633 2 MOAI1S $T=806620 799800 1 0 $X=806620 $Y=794380
X3865 4505 926 1 4505 4361 4652 2 MOAI1S $T=807860 819960 0 0 $X=807860 $Y=819580
X3866 4544 4647 1 4544 848 4653 2 MOAI1S $T=809720 890520 1 0 $X=809720 $Y=885100
X3867 4645 930 1 4645 881 4661 2 MOAI1S $T=810340 739320 1 0 $X=810340 $Y=733900
X3868 4702 4658 1 4702 4646 4641 2 MOAI1S $T=823360 870360 0 180 $X=819640 $Y=864940
X3869 4702 944 1 4702 4437 4663 2 MOAI1S $T=823980 850200 1 180 $X=820260 $Y=849820
X3870 947 4708 1 904 941 4698 2 MOAI1S $T=825220 900600 0 180 $X=821500 $Y=895180
X3871 4731 4703 1 4731 4437 4727 2 MOAI1S $T=827700 860280 0 180 $X=823980 $Y=854860
X3872 4716 954 1 4716 4590 4697 2 MOAI1S $T=834520 890520 0 180 $X=830800 $Y=885100
X3873 4539 4771 1 4539 551 4784 2 MOAI1S $T=831420 789720 1 0 $X=831420 $Y=784300
X3874 4788 4792 1 4788 4646 4797 2 MOAI1S $T=833900 870360 1 0 $X=833900 $Y=864940
X3875 4788 4563 1 4788 4590 4804 2 MOAI1S $T=833900 880440 1 0 $X=833900 $Y=875020
X3876 4716 4781 1 4716 4815 4807 2 MOAI1S $T=837620 890520 0 0 $X=837620 $Y=890140
X3877 4840 4625 1 4840 4590 4838 2 MOAI1S $T=847540 880440 1 180 $X=843820 $Y=880060
X3878 4788 4846 1 4788 4815 4832 2 MOAI1S $T=845060 890520 0 0 $X=845060 $Y=890140
X3879 4840 4336 1 4840 4710 4869 2 MOAI1S $T=846920 880440 1 0 $X=846920 $Y=875020
X3880 4840 4870 1 4840 4815 4860 2 MOAI1S $T=851260 880440 1 180 $X=847540 $Y=880060
X3881 4822 4502 1 4822 4646 4877 2 MOAI1S $T=848160 870360 1 0 $X=848160 $Y=864940
X3882 4814 4751 1 4814 4646 4873 2 MOAI1S $T=848780 860280 1 0 $X=848780 $Y=854860
X3883 4882 4889 1 4882 978 4913 2 MOAI1S $T=852500 880440 0 0 $X=852500 $Y=880060
X3884 4882 979 1 4882 4710 4937 2 MOAI1S $T=858700 880440 1 0 $X=858700 $Y=875020
X3885 5427 5439 1 5427 5435 5404 2 MOAI1S $T=954180 779640 0 180 $X=950460 $Y=774220
X3886 5379 1076 1 5379 5435 5466 2 MOAI1S $T=952320 789720 0 0 $X=952320 $Y=789340
X3887 5325 5504 1 5325 5496 5492 2 MOAI1S $T=964100 880440 0 180 $X=960380 $Y=875020
X3888 5427 5500 1 5427 5496 5507 2 MOAI1S $T=961620 779640 0 0 $X=961620 $Y=779260
X3889 5330 5478 1 5330 5496 5517 2 MOAI1S $T=962240 789720 1 0 $X=962240 $Y=784300
X3890 5379 5508 1 5379 5496 5516 2 MOAI1S $T=964100 799800 1 0 $X=964100 $Y=794380
X3891 5304 5510 1 5304 5496 5519 2 MOAI1S $T=964100 860280 0 0 $X=964100 $Y=859900
X3892 5345 5522 1 5345 5496 5509 2 MOAI1S $T=968440 809880 1 180 $X=964720 $Y=809500
X3893 5653 5654 1 5653 1110 5627 2 MOAI1S $T=991380 809880 0 0 $X=991380 $Y=809500
X3894 5659 5668 1 5659 1110 5622 2 MOAI1S $T=996960 860280 0 180 $X=993240 $Y=854860
X3895 5665 5670 1 5665 1110 5635 2 MOAI1S $T=997580 789720 1 180 $X=993860 $Y=789340
X3896 5666 5669 1 5666 1115 5676 2 MOAI1S $T=995100 890520 1 0 $X=995100 $Y=885100
X3897 5671 5683 1 5671 1110 5628 2 MOAI1S $T=999440 809880 1 180 $X=995720 $Y=809500
X3898 5659 5695 1 5659 1115 5664 2 MOAI1S $T=1000680 860280 1 180 $X=996960 $Y=859900
X3899 5677 5672 1 5677 1114 5699 2 MOAI1S $T=997580 739320 1 0 $X=997580 $Y=733900
X3900 1118 1120 1 1118 1114 1116 2 MOAI1S $T=1002540 729240 0 180 $X=998820 $Y=723820
X3901 5698 1123 1 5698 1115 5631 2 MOAI1S $T=1003160 900600 0 180 $X=999440 $Y=895180
X3902 5714 5727 1 5714 1122 5696 2 MOAI1S $T=1004400 880440 0 180 $X=1000680 $Y=875020
X3903 5653 1126 1 5653 5745 5713 2 MOAI1S $T=1003160 809880 0 0 $X=1003160 $Y=809500
X3904 5733 5762 1 5733 5745 5743 2 MOAI1S $T=1009360 789720 1 180 $X=1005640 $Y=789340
X3905 5735 1130 1 5735 1115 5753 2 MOAI1S $T=1005640 860280 1 0 $X=1005640 $Y=854860
X3906 5720 5731 1 5720 5745 5792 2 MOAI1S $T=1006260 779640 1 0 $X=1006260 $Y=774220
X3907 5736 5770 1 5736 1134 5751 2 MOAI1S $T=1010600 739320 1 180 $X=1006880 $Y=738940
X3908 5773 5697 1 5697 5760 5710 2 MOAI1S $T=1010600 840120 0 180 $X=1006880 $Y=834700
X3909 5671 5772 1 5671 5745 5721 2 MOAI1S $T=1011220 799800 1 180 $X=1007500 $Y=799420
X3910 5724 1137 1 5724 5755 5738 2 MOAI1S $T=1012460 880440 1 180 $X=1008740 $Y=880060
X3911 5665 5785 1 5665 5745 5769 2 MOAI1S $T=1013700 789720 1 180 $X=1009980 $Y=789340
X3912 5775 1136 1 5775 1122 5788 2 MOAI1S $T=1009980 880440 1 0 $X=1009980 $Y=875020
X3913 5781 5799 1 5781 1144 5787 2 MOAI1S $T=1016800 850200 0 180 $X=1013080 $Y=844780
X3914 5724 5791 1 5724 5501 5811 2 MOAI1S $T=1013080 890520 0 0 $X=1013080 $Y=890140
X3915 5796 5804 1 5796 1134 5722 2 MOAI1S $T=1018040 749400 0 180 $X=1014320 $Y=743980
X3916 5794 5771 1 5794 1144 5783 2 MOAI1S $T=1018040 860280 1 180 $X=1014320 $Y=859900
X3917 5796 5815 1 5796 1147 5780 2 MOAI1S $T=1019280 759480 0 180 $X=1015560 $Y=754060
X3918 5797 5801 1 5797 5760 5718 2 MOAI1S $T=1015560 830040 1 0 $X=1015560 $Y=824620
X3919 5775 5807 1 5775 1149 1151 2 MOAI1S $T=1016180 900600 1 0 $X=1016180 $Y=895180
X3920 5802 5702 1 5802 5501 5810 2 MOAI1S $T=1020520 850200 0 180 $X=1016800 $Y=844780
X3921 5775 5688 1 5775 1144 5824 2 MOAI1S $T=1017420 880440 1 0 $X=1017420 $Y=875020
X3922 5736 5816 1 5736 1147 5825 2 MOAI1S $T=1018040 739320 0 0 $X=1018040 $Y=738940
X3923 5701 5823 1 5701 5817 5795 2 MOAI1S $T=1021760 809880 0 180 $X=1018040 $Y=804460
X3924 5797 5827 1 5797 5501 5818 2 MOAI1S $T=1023000 830040 0 180 $X=1019280 $Y=824620
X3925 5733 5833 1 5733 5435 5809 2 MOAI1S $T=1023620 779640 1 180 $X=1019900 $Y=779260
X3926 5826 5834 1 5826 5760 5814 2 MOAI1S $T=1023620 819960 0 180 $X=1019900 $Y=814540
X3927 5830 1157 1 5830 1147 5808 2 MOAI1S $T=1024860 729240 0 180 $X=1021140 $Y=723820
X3928 5720 5843 1 5720 5435 5813 2 MOAI1S $T=1025480 759480 0 180 $X=1021760 $Y=754060
X3929 5870 5871 1 5870 5817 5793 2 MOAI1S $T=1031060 799800 0 180 $X=1027340 $Y=794380
X3930 5863 5899 1 5863 5887 5837 2 MOAI1S $T=1034160 759480 0 180 $X=1030440 $Y=754060
X3931 1166 5903 1 1166 5755 5883 2 MOAI1S $T=1034160 880440 1 180 $X=1030440 $Y=880060
X3932 5888 5908 1 5888 5887 5867 2 MOAI1S $T=1034780 779640 1 180 $X=1031060 $Y=779260
X3933 5826 5892 1 5826 5890 5919 2 MOAI1S $T=1031060 819960 0 0 $X=1031060 $Y=819580
X3934 5803 5915 1 5803 1170 5894 2 MOAI1S $T=1036020 739320 0 180 $X=1032300 $Y=733900
X3935 5922 5902 1 5902 5760 5901 2 MOAI1S $T=1036640 850200 0 180 $X=1032920 $Y=844780
X3936 1166 1174 1 1166 1149 5905 2 MOAI1S $T=1036640 900600 0 180 $X=1032920 $Y=895180
X3937 5796 5916 1 5878 5887 5932 2 MOAI1S $T=1034160 759480 1 0 $X=1034160 $Y=754060
X3938 1166 5917 1 5923 1144 5822 2 MOAI1S $T=1034160 860280 0 0 $X=1034160 $Y=859900
X3939 1162 5886 1 1162 1170 1172 2 MOAI1S $T=1039120 729240 0 180 $X=1035400 $Y=723820
X3940 5900 5927 1 5900 5887 5942 2 MOAI1S $T=1036020 809880 0 0 $X=1036020 $Y=809500
X3941 5923 5937 1 5923 5760 5906 2 MOAI1S $T=1040360 850200 0 180 $X=1036640 $Y=844780
X3942 5878 5945 1 5878 5939 5893 2 MOAI1S $T=1041600 759480 0 180 $X=1037880 $Y=754060
X3943 5926 5950 1 5926 1144 5913 2 MOAI1S $T=1042220 860280 1 180 $X=1038500 $Y=859900
X3944 1177 5951 1 1177 5755 5938 2 MOAI1S $T=1042220 890520 0 180 $X=1038500 $Y=885100
X3945 5955 5976 1 5955 5935 5947 2 MOAI1S $T=1046560 809880 1 180 $X=1042840 $Y=809500
X3946 5803 5969 1 5803 1168 5983 2 MOAI1S $T=1044080 739320 0 0 $X=1044080 $Y=738940
X3947 5863 1186 1 5863 5939 5995 2 MOAI1S $T=1046560 759480 1 0 $X=1046560 $Y=754060
X3948 5900 5992 1 5900 5935 6010 2 MOAI1S $T=1048420 799800 0 0 $X=1048420 $Y=799420
X3949 5888 6001 1 5888 5935 6013 2 MOAI1S $T=1049660 779640 0 0 $X=1049660 $Y=779260
X3950 5910 6002 1 5910 5935 5989 2 MOAI1S $T=1049660 789720 0 0 $X=1049660 $Y=789340
X3951 1367 2 1336 1340 1 NR2 $T=228780 830040 0 0 $X=228780 $Y=829660
X3952 15 2 1344 1384 1 NR2 $T=233120 789720 0 180 $X=231260 $Y=784300
X3953 1397 2 1364 1352 1 NR2 $T=233120 850200 1 180 $X=231260 $Y=849820
X3954 1373 2 1379 1409 1 NR2 $T=231880 819960 0 0 $X=231880 $Y=819580
X3955 1390 2 1426 1396 1 NR2 $T=231880 830040 0 0 $X=231880 $Y=829660
X3956 1390 2 1424 1409 1 NR2 $T=231880 840120 1 0 $X=231880 $Y=834700
X3957 15 2 1415 1396 1 NR2 $T=234360 830040 0 180 $X=232500 $Y=824620
X3958 1373 2 1392 1408 1 NR2 $T=233120 769560 1 0 $X=233120 $Y=764140
X3959 1373 2 1387 1412 1 NR2 $T=233120 779640 0 0 $X=233120 $Y=779260
X3960 1390 2 1405 1384 1 NR2 $T=234980 789720 0 180 $X=233120 $Y=784300
X3961 1400 2 1383 1409 1 NR2 $T=233120 799800 1 0 $X=233120 $Y=794380
X3962 1407 2 1378 1418 1 NR2 $T=233740 759480 0 0 $X=233740 $Y=759100
X3963 15 2 1385 1412 1 NR2 $T=233740 799800 0 0 $X=233740 $Y=799420
X3964 1407 2 1406 1409 1 NR2 $T=235600 809880 1 180 $X=233740 $Y=809500
X3965 1407 2 1393 1411 1 NR2 $T=236220 779640 0 180 $X=234360 $Y=774220
X3966 1373 2 1425 1411 1 NR2 $T=234360 819960 1 0 $X=234360 $Y=814540
X3967 15 2 1389 1411 1 NR2 $T=234980 819960 0 0 $X=234980 $Y=819580
X3968 1400 2 1388 1421 1 NR2 $T=237460 759480 1 180 $X=235600 $Y=759100
X3969 1400 2 1422 1433 1 NR2 $T=235600 799800 1 0 $X=235600 $Y=794380
X3970 1400 2 1410 1396 1 NR2 $T=236840 789720 1 0 $X=236840 $Y=784300
X3971 1390 2 1427 1412 1 NR2 $T=238700 799800 1 180 $X=236840 $Y=799420
X3972 1390 2 1434 1411 1 NR2 $T=239940 819960 1 180 $X=238080 $Y=819580
X3973 1407 2 1440 1408 1 NR2 $T=240560 779640 0 180 $X=238700 $Y=774220
X3974 1390 2 1445 1433 1 NR2 $T=238700 830040 0 0 $X=238700 $Y=829660
X3975 15 2 1431 1409 1 NR2 $T=240560 840120 0 180 $X=238700 $Y=834700
X3976 15 2 1449 1433 1 NR2 $T=241180 830040 0 0 $X=241180 $Y=829660
X3977 1407 2 1466 1396 1 NR2 $T=242420 799800 0 0 $X=242420 $Y=799420
X3978 1493 2 1491 1396 1 NR2 $T=245520 779640 1 180 $X=243660 $Y=779260
X3979 1407 2 1488 1433 1 NR2 $T=244280 819960 0 0 $X=244280 $Y=819580
X3980 1493 2 1476 1433 1 NR2 $T=247380 799800 1 180 $X=245520 $Y=799420
X3981 36 2 1506 1500 1 NR2 $T=248000 749400 1 0 $X=248000 $Y=743980
X3982 1493 2 1513 1408 1 NR2 $T=249240 749400 0 0 $X=249240 $Y=749020
X3983 44 2 1501 1421 1 NR2 $T=251100 759480 0 180 $X=249240 $Y=754060
X3984 1545 2 40 46 1 NR2 $T=252960 900600 0 180 $X=251100 $Y=895180
X3985 1347 2 1530 1525 1 NR2 $T=252960 809880 0 0 $X=252960 $Y=809500
X3986 29 2 1538 1532 1 NR2 $T=254820 779640 0 0 $X=254820 $Y=779260
X3987 50 2 1526 1532 1 NR2 $T=255440 749400 0 0 $X=255440 $Y=749020
X3988 56 2 1546 1568 1 NR2 $T=258540 880440 1 0 $X=258540 $Y=875020
X3989 1581 2 1484 1547 1 NR2 $T=261640 759480 0 180 $X=259780 $Y=754060
X3990 1518 2 1576 1485 1 NR2 $T=259780 809880 1 0 $X=259780 $Y=804460
X3991 1514 2 1565 1563 1 NR2 $T=259780 819960 1 0 $X=259780 $Y=814540
X3992 50 2 1566 1408 1 NR2 $T=261640 759480 0 0 $X=261640 $Y=759100
X3993 1493 2 1590 1409 1 NR2 $T=261640 789720 0 0 $X=261640 $Y=789340
X3994 63 2 1505 1568 1 NR2 $T=263500 880440 1 180 $X=261640 $Y=880060
X3995 50 2 1569 1500 1 NR2 $T=263500 739320 0 0 $X=263500 $Y=738940
X3996 67 2 1582 1532 1 NR2 $T=265360 789720 0 180 $X=263500 $Y=784300
X3997 1595 2 1535 65 1 NR2 $T=265980 890520 0 180 $X=264120 $Y=885100
X3998 1581 2 1575 1421 1 NR2 $T=265360 759480 0 0 $X=265360 $Y=759100
X3999 1581 2 1605 1418 1 NR2 $T=267220 739320 0 0 $X=267220 $Y=738940
X4000 20 2 1614 1622 1 NR2 $T=267220 749400 1 0 $X=267220 $Y=743980
X4001 67 2 1603 1500 1 NR2 $T=267220 779640 1 0 $X=267220 $Y=774220
X4002 1565 2 1606 1576 1 NR2 $T=269080 799800 1 180 $X=267220 $Y=799420
X4003 29 2 1611 1500 1 NR2 $T=268460 759480 0 0 $X=268460 $Y=759100
X4004 1568 2 1623 1549 1 NR2 $T=270320 870360 1 0 $X=270320 $Y=864940
X4005 1493 2 1629 1418 1 NR2 $T=272800 759480 0 180 $X=270940 $Y=754060
X4006 1581 2 1617 1638 1 NR2 $T=270940 779640 0 0 $X=270940 $Y=779260
X4007 1644 2 1639 1421 1 NR2 $T=275900 739320 0 180 $X=274040 $Y=733900
X4008 1644 2 1633 1638 1 NR2 $T=275900 779640 1 180 $X=274040 $Y=779260
X4009 29 2 1664 1622 1 NR2 $T=275900 769560 1 0 $X=275900 $Y=764140
X4010 1644 2 1656 1547 1 NR2 $T=275900 769560 0 0 $X=275900 $Y=769180
X4011 1493 2 1665 1532 1 NR2 $T=277760 749400 0 0 $X=277760 $Y=749020
X4012 36 2 1637 1532 1 NR2 $T=277760 759480 1 0 $X=277760 $Y=754060
X4013 71 2 1627 87 1 NR2 $T=277760 870360 0 0 $X=277760 $Y=869980
X4014 1644 2 1673 1418 1 NR2 $T=280240 739320 0 180 $X=278380 $Y=733900
X4015 67 2 1689 1622 1 NR2 $T=279620 769560 0 0 $X=279620 $Y=769180
X4016 1581 2 1683 1408 1 NR2 $T=281480 759480 1 0 $X=281480 $Y=754060
X4017 1549 2 1679 87 1 NR2 $T=283340 860280 1 180 $X=281480 $Y=859900
X4018 71 2 1686 91 1 NR2 $T=281480 870360 1 0 $X=281480 $Y=864940
X4019 36 2 1700 1622 1 NR2 $T=284580 749400 0 180 $X=282720 $Y=743980
X4020 20 2 1684 1500 1 NR2 $T=285200 759480 0 180 $X=283340 $Y=754060
X4021 1685 2 1680 91 1 NR2 $T=287060 890520 0 180 $X=285200 $Y=885100
X4022 95 2 1697 1685 1 NR2 $T=285200 890520 0 0 $X=285200 $Y=890140
X4023 1751 2 1730 1704 1 NR2 $T=288300 779640 0 180 $X=286440 $Y=774220
X4024 1738 2 1725 100 1 NR2 $T=292020 890520 0 180 $X=290160 $Y=885100
X4025 20 2 1710 1740 1 NR2 $T=290780 749400 1 0 $X=290780 $Y=743980
X4026 1751 2 1766 1421 1 NR2 $T=293880 739320 0 0 $X=293880 $Y=738940
X4027 1751 2 1776 1547 1 NR2 $T=293880 769560 1 0 $X=293880 $Y=764140
X4028 1751 2 1736 1638 1 NR2 $T=293880 779640 1 0 $X=293880 $Y=774220
X4029 1777 2 1749 1752 1 NR2 $T=295740 870360 1 180 $X=293880 $Y=869980
X4030 107 2 1729 100 1 NR2 $T=295740 900600 0 180 $X=293880 $Y=895180
X4031 29 2 1784 1740 1 NR2 $T=295120 769560 0 0 $X=295120 $Y=769180
X4032 1772 2 1759 1752 1 NR2 $T=296980 880440 1 180 $X=295120 $Y=880060
X4033 1773 2 1737 112 1 NR2 $T=296360 890520 0 0 $X=296360 $Y=890140
X4034 107 2 1771 1777 1 NR2 $T=297600 880440 0 0 $X=297600 $Y=880060
X4035 114 2 1761 111 1 NR2 $T=299460 900600 0 180 $X=297600 $Y=895180
X4036 67 2 1778 1740 1 NR2 $T=298840 779640 1 0 $X=298840 $Y=774220
X4037 117 2 1743 116 1 NR2 $T=302560 900600 0 180 $X=300700 $Y=895180
X4038 1773 2 119 121 1 NR2 $T=301940 890520 0 0 $X=301940 $Y=890140
X4039 116 2 1806 122 1 NR2 $T=302560 900600 1 0 $X=302560 $Y=895180
X4040 1773 2 1838 129 1 NR2 $T=310000 870360 0 0 $X=310000 $Y=869980
X4041 143 2 1862 1704 1 NR2 $T=313720 779640 1 180 $X=311860 $Y=779260
X4042 1861 2 1647 129 1 NR2 $T=313720 870360 1 180 $X=311860 $Y=869980
X4043 1861 2 1840 1857 1 NR2 $T=313720 880440 0 180 $X=311860 $Y=875020
X4044 136 2 140 129 1 NR2 $T=313720 900600 0 180 $X=311860 $Y=895180
X4045 1869 2 1839 135 1 NR2 $T=314960 880440 1 180 $X=313100 $Y=880060
X4046 135 2 1836 1871 1 NR2 $T=313720 890520 1 0 $X=313720 $Y=885100
X4047 151 2 1845 1871 1 NR2 $T=316820 870360 0 180 $X=314960 $Y=864940
X4048 1869 2 147 146 1 NR2 $T=314960 890520 0 0 $X=314960 $Y=890140
X4049 97 2 1859 1704 1 NR2 $T=319920 789720 0 180 $X=318060 $Y=784300
X4050 67 2 1889 1885 1 NR2 $T=318680 779640 0 0 $X=318680 $Y=779260
X4051 67 2 1879 1955 1 NR2 $T=319920 789720 1 0 $X=319920 $Y=784300
X4052 146 2 1894 1772 1 NR2 $T=322400 890520 1 180 $X=320540 $Y=890140
X4053 110 2 1910 1547 1 NR2 $T=323640 769560 0 0 $X=323640 $Y=769180
X4054 165 2 1950 164 1 NR2 $T=327360 880440 0 0 $X=327360 $Y=880060
X4055 167 2 1953 136 1 NR2 $T=327980 890520 0 0 $X=327980 $Y=890140
X4056 172 2 1904 136 1 NR2 $T=331080 870360 1 180 $X=329220 $Y=869980
X4057 60 2 1954 1861 1 NR2 $T=330460 880440 0 0 $X=330460 $Y=880060
X4058 61 2 182 1773 1 NR2 $T=336660 880440 1 180 $X=334800 $Y=880060
X4059 183 2 1990 2020 1 NR2 $T=337900 799800 1 0 $X=337900 $Y=794380
X4060 1954 2 2035 182 1 NR2 $T=338520 880440 0 0 $X=338520 $Y=880060
X4061 158 2 191 193 1 NR2 $T=339760 900600 1 0 $X=339760 $Y=895180
X4062 2045 2 192 2035 1 NR2 $T=342860 880440 1 180 $X=341000 $Y=880060
X4063 151 2 1914 2065 1 NR2 $T=344720 880440 1 0 $X=344720 $Y=875020
X4064 2084 2 2092 202 1 NR2 $T=348440 759480 0 0 $X=348440 $Y=759100
X4065 2084 2 2075 199 1 NR2 $T=350300 779640 1 180 $X=348440 $Y=779260
X4066 2113 2 2088 199 1 NR2 $T=350920 769560 1 180 $X=349060 $Y=769180
X4067 2084 2 2094 2125 1 NR2 $T=350920 779640 1 0 $X=350920 $Y=774220
X4068 2084 2 1797 2121 1 NR2 $T=350920 779640 0 0 $X=350920 $Y=779260
X4069 2113 2 2116 202 1 NR2 $T=352160 759480 1 0 $X=352160 $Y=754060
X4070 2113 2 2040 2121 1 NR2 $T=352160 769560 0 0 $X=352160 $Y=769180
X4071 2168 2 2128 202 1 NR2 $T=357740 729240 1 180 $X=355880 $Y=728860
X4072 205 2 2124 212 1 NR2 $T=355880 739320 0 0 $X=355880 $Y=738940
X4073 2084 2 2062 2150 1 NR2 $T=355880 779640 0 0 $X=355880 $Y=779260
X4074 164 2 2143 1911 1 NR2 $T=357740 880440 0 180 $X=355880 $Y=875020
X4075 213 2 2130 207 1 NR2 $T=359600 739320 0 180 $X=357740 $Y=733900
X4076 2113 2 2179 212 1 NR2 $T=359600 739320 0 0 $X=359600 $Y=738940
X4077 2168 2 2167 2121 1 NR2 $T=363940 769560 1 180 $X=362080 $Y=769180
X4078 2168 2 2176 199 1 NR2 $T=364560 759480 1 180 $X=362700 $Y=759100
X4079 2184 2 2178 202 1 NR2 $T=365180 729240 1 180 $X=363320 $Y=728860
X4080 2168 2 2137 211 1 NR2 $T=364560 759480 0 0 $X=364560 $Y=759100
X4081 2151 2 2204 226 1 NR2 $T=364560 809880 0 0 $X=364560 $Y=809500
X4082 129 2 2162 2100 1 NR2 $T=364560 890520 1 0 $X=364560 $Y=885100
X4083 213 2 228 212 1 NR2 $T=368280 729240 0 180 $X=366420 $Y=723820
X4084 2184 2 2192 199 1 NR2 $T=368280 759480 0 180 $X=366420 $Y=754060
X4085 1912 2 2205 2100 1 NR2 $T=368280 890520 0 180 $X=366420 $Y=885100
X4086 2168 2 2201 2125 1 NR2 $T=367040 759480 0 0 $X=367040 $Y=759100
X4087 2209 2 2202 2125 1 NR2 $T=368900 779640 1 180 $X=367040 $Y=779260
X4088 229 2 2166 233 1 NR2 $T=367040 890520 0 0 $X=367040 $Y=890140
X4089 1869 2 2198 236 1 NR2 $T=368280 900600 1 0 $X=368280 $Y=895180
X4090 2184 2 2267 2150 1 NR2 $T=370140 759480 1 0 $X=370140 $Y=754060
X4091 2184 2 2207 2121 1 NR2 $T=370140 759480 0 0 $X=370140 $Y=759100
X4092 2209 2 2187 2150 1 NR2 $T=370140 789720 1 0 $X=370140 $Y=784300
X4093 158 2 2241 101 1 NR2 $T=370140 890520 0 0 $X=370140 $Y=890140
X4094 2065 2 2230 2236 1 NR2 $T=371380 870360 1 0 $X=371380 $Y=864940
X4095 2168 2 2228 2150 1 NR2 $T=373860 779640 0 180 $X=372000 $Y=774220
X4096 1869 2 239 238 1 NR2 $T=372000 900600 1 0 $X=372000 $Y=895180
X4097 245 2 2252 242 1 NR2 $T=376340 799800 0 180 $X=374480 $Y=794380
X4098 203 2 2254 100 1 NR2 $T=374480 890520 1 0 $X=374480 $Y=885100
X4099 2255 2 244 202 1 NR2 $T=375100 729240 1 0 $X=375100 $Y=723820
X4100 2255 2 2239 199 1 NR2 $T=375100 739320 0 0 $X=375100 $Y=738940
X4101 2184 2 2249 211 1 NR2 $T=375100 749400 1 0 $X=375100 $Y=743980
X4102 2204 2 2262 2263 1 NR2 $T=375100 809880 1 0 $X=375100 $Y=804460
X4103 2250 2 2263 157 1 NR2 $T=375720 819960 1 0 $X=375720 $Y=814540
X4104 1871 2 2270 236 1 NR2 $T=375720 880440 1 0 $X=375720 $Y=875020
X4105 1871 2 2258 2236 1 NR2 $T=377580 880440 1 180 $X=375720 $Y=880060
X4106 2184 2 2259 2125 1 NR2 $T=376340 749400 0 0 $X=376340 $Y=749020
X4107 247 2 2265 101 1 NR2 $T=378200 890520 0 180 $X=376340 $Y=885100
X4108 247 2 2274 100 1 NR2 $T=376960 900600 1 0 $X=376960 $Y=895180
X4109 235 2 2261 2061 1 NR2 $T=377580 880440 0 0 $X=377580 $Y=880060
X4110 249 2 2272 2061 1 NR2 $T=378200 890520 1 0 $X=378200 $Y=885100
X4111 2255 2 2297 2150 1 NR2 $T=378820 749400 0 0 $X=378820 $Y=749020
X4112 2255 2 2256 2121 1 NR2 $T=378820 759480 1 0 $X=378820 $Y=754060
X4113 172 2 2279 2300 1 NR2 $T=378820 880440 1 0 $X=378820 $Y=875020
X4114 257 2 2286 199 1 NR2 $T=384400 729240 0 180 $X=382540 $Y=723820
X4115 257 2 2331 254 1 NR2 $T=386260 739320 0 180 $X=384400 $Y=733900
X4116 257 2 2345 2125 1 NR2 $T=386260 729240 1 0 $X=386260 $Y=723820
X4117 257 2 2346 2150 1 NR2 $T=386260 739320 1 0 $X=386260 $Y=733900
X4118 188 2 2313 259 1 NR2 $T=386260 890520 1 0 $X=386260 $Y=885100
X4119 2177 2 2322 253 1 NR2 $T=388120 799800 0 0 $X=388120 $Y=799420
X4120 261 2 267 265 1 NR2 $T=389980 729240 1 0 $X=389980 $Y=723820
X4121 261 2 2361 2121 1 NR2 $T=391840 739320 0 180 $X=389980 $Y=733900
X4122 1886 2 2367 218 1 NR2 $T=393080 840120 0 180 $X=391220 $Y=834700
X4123 2310 2 2074 269 1 NR2 $T=391220 890520 0 0 $X=391220 $Y=890140
X4124 2376 2 2302 2322 1 NR2 $T=393700 809880 0 180 $X=391840 $Y=804460
X4125 1912 2 2445 2061 1 NR2 $T=394940 890520 1 0 $X=394940 $Y=885100
X4126 2400 2 2376 273 1 NR2 $T=398040 799800 1 180 $X=396180 $Y=799420
X4127 2425 2 2409 2404 1 NR2 $T=400520 850200 0 180 $X=398660 $Y=844780
X4128 2330 2 2404 177 1 NR2 $T=398660 860280 1 0 $X=398660 $Y=854860
X4129 280 2 281 2300 1 NR2 $T=399900 900600 1 0 $X=399900 $Y=895180
X4130 235 2 282 2300 1 NR2 $T=400520 890520 0 0 $X=400520 $Y=890140
X4131 270 2 283 252 1 NR2 $T=403620 900600 0 180 $X=401760 $Y=895180
X4132 2451 2 2426 2438 1 NR2 $T=405480 779640 0 180 $X=403620 $Y=774220
X4133 2456 2 2432 2438 1 NR2 $T=406100 789720 0 180 $X=404240 $Y=784300
X4134 2397 2 2425 171 1 NR2 $T=406100 840120 1 180 $X=404240 $Y=839740
X4135 288 2 2428 2438 1 NR2 $T=407340 749400 1 180 $X=405480 $Y=749020
X4136 2456 2 2449 286 1 NR2 $T=405480 759480 0 0 $X=405480 $Y=759100
X4137 2465 2 2457 285 1 NR2 $T=407340 769560 1 180 $X=405480 $Y=769180
X4138 2451 2 2454 286 1 NR2 $T=406100 759480 1 0 $X=406100 $Y=754060
X4139 2468 2 2443 286 1 NR2 $T=407960 779640 0 180 $X=406100 $Y=774220
X4140 288 2 2448 2474 1 NR2 $T=407340 749400 1 0 $X=407340 $Y=743980
X4141 2465 2 2464 286 1 NR2 $T=409200 789720 0 180 $X=407340 $Y=784300
X4142 2476 2 2444 1969 1 NR2 $T=409200 830040 0 180 $X=407340 $Y=824620
X4143 270 2 2479 290 1 NR2 $T=407340 900600 1 0 $X=407340 $Y=895180
X4144 2468 2 2455 285 1 NR2 $T=409820 769560 0 180 $X=407960 $Y=764140
X4145 2468 2 2486 2489 1 NR2 $T=407960 769560 0 0 $X=407960 $Y=769180
X4146 2465 2 2466 293 1 NR2 $T=409200 779640 1 0 $X=409200 $Y=774220
X4147 2465 2 2480 2438 1 NR2 $T=409200 789720 1 0 $X=409200 $Y=784300
X4148 2209 2 2485 2438 1 NR2 $T=409200 799800 1 0 $X=409200 $Y=794380
X4149 295 2 2495 2438 1 NR2 $T=412920 729240 1 180 $X=411060 $Y=728860
X4150 2465 2 2424 296 1 NR2 $T=411060 759480 0 0 $X=411060 $Y=759100
X4151 2465 2 2498 2474 1 NR2 $T=411680 789720 1 0 $X=411680 $Y=784300
X4152 2451 2 2501 2474 1 NR2 $T=414160 769560 1 180 $X=412300 $Y=769180
X4153 2209 2 2504 2474 1 NR2 $T=412920 799800 1 0 $X=412920 $Y=794380
X4154 2209 2 2511 293 1 NR2 $T=414160 789720 1 0 $X=414160 $Y=784300
X4155 2451 2 2526 293 1 NR2 $T=414780 769560 0 0 $X=414780 $Y=769180
X4156 2456 2 2531 2489 1 NR2 $T=416020 779640 0 0 $X=416020 $Y=779260
X4157 2456 2 2535 2474 1 NR2 $T=416020 789720 0 0 $X=416020 $Y=789340
X4158 2451 2 2534 2489 1 NR2 $T=417880 769560 0 0 $X=417880 $Y=769180
X4159 295 2 2524 293 1 NR2 $T=418500 739320 0 0 $X=418500 $Y=738940
X4160 295 2 2503 2489 1 NR2 $T=418500 749400 0 0 $X=418500 $Y=749020
X4161 295 2 2544 285 1 NR2 $T=419740 729240 1 0 $X=419740 $Y=723820
X4162 288 2 2539 2489 1 NR2 $T=421600 759480 0 180 $X=419740 $Y=754060
X4163 288 2 2556 285 1 NR2 $T=421600 739320 0 0 $X=421600 $Y=738940
X4164 287 2 2563 291 1 NR2 $T=422840 729240 1 0 $X=422840 $Y=723820
X4165 2413 2 2569 296 1 NR2 $T=423460 749400 0 0 $X=423460 $Y=749020
X4166 2413 2 2568 294 1 NR2 $T=425320 739320 0 0 $X=425320 $Y=738940
X4167 301 2 2577 285 1 NR2 $T=425320 759480 1 0 $X=425320 $Y=754060
X4168 2468 2 2557 296 1 NR2 $T=427180 769560 0 180 $X=425320 $Y=764140
X4169 2456 2 2566 285 1 NR2 $T=426560 759480 0 0 $X=426560 $Y=759100
X4170 2456 2 2564 293 1 NR2 $T=426560 779640 1 0 $X=426560 $Y=774220
X4171 298 2 2646 333 1 NR2 $T=439580 749400 1 0 $X=439580 $Y=743980
X4172 292 2 2647 333 1 NR2 $T=439580 749400 0 0 $X=439580 $Y=749020
X4173 298 2 2654 339 1 NR2 $T=441440 739320 0 0 $X=441440 $Y=738940
X4174 292 2 2673 342 1 NR2 $T=446400 729240 1 0 $X=446400 $Y=723820
X4175 2413 2 2663 333 1 NR2 $T=446400 739320 1 0 $X=446400 $Y=733900
X4176 2413 2 2711 339 1 NR2 $T=451980 729240 0 0 $X=451980 $Y=728860
X4177 358 2 2714 339 1 NR2 $T=456940 729240 1 180 $X=455080 $Y=728860
X4178 379 2 2839 2819 1 NR2 $T=476780 729240 0 180 $X=474920 $Y=723820
X4179 3165 2 3168 452 1 NR2 $T=537540 850200 0 0 $X=537540 $Y=849820
X4180 3173 2 3169 454 1 NR2 $T=540640 880440 1 0 $X=540640 $Y=875020
X4181 461 2 3197 3120 1 NR2 $T=544360 890520 0 180 $X=542500 $Y=885100
X4182 460 2 3187 3208 1 NR2 $T=546220 809880 0 0 $X=546220 $Y=809500
X4183 3234 2 3181 475 1 NR2 $T=554900 789720 0 0 $X=554900 $Y=789340
X4184 3296 2 3319 3138 1 NR2 $T=566680 799800 1 0 $X=566680 $Y=794380
X4185 3333 2 3321 454 1 NR2 $T=571020 870360 0 180 $X=569160 $Y=864940
X4186 3414 2 3417 475 1 NR2 $T=583420 789720 1 0 $X=583420 $Y=784300
X4187 3480 2 3137 3491 1 NR2 $T=597680 789720 1 0 $X=597680 $Y=784300
X4188 546 2 3404 3486 1 NR2 $T=602020 789720 1 180 $X=600160 $Y=789340
X4189 3507 2 494 3486 1 NR2 $T=602640 789720 0 180 $X=600780 $Y=784300
X4190 3173 2 3494 520 1 NR2 $T=602640 880440 0 180 $X=600780 $Y=875020
X4191 3507 2 3495 3491 1 NR2 $T=603260 779640 1 180 $X=601400 $Y=779260
X4192 3532 2 3315 3491 1 NR2 $T=606360 779640 1 180 $X=604500 $Y=779260
X4193 3532 2 3472 3486 1 NR2 $T=608840 779640 0 180 $X=606980 $Y=774220
X4194 3596 2 3601 3613 1 NR2 $T=620620 809880 1 0 $X=620620 $Y=804460
X4195 3611 2 3629 3436 1 NR2 $T=624340 779640 1 0 $X=624340 $Y=774220
X4196 3333 2 3627 593 1 NR2 $T=624340 880440 1 0 $X=624340 $Y=875020
X4197 3173 2 3656 593 1 NR2 $T=629920 880440 1 0 $X=629920 $Y=875020
X4198 3234 2 3707 603 1 NR2 $T=641080 799800 1 0 $X=641080 $Y=794380
X4199 3414 2 3607 603 1 NR2 $T=641700 769560 0 0 $X=641700 $Y=769180
X4200 546 2 3761 3491 1 NR2 $T=656580 779640 0 0 $X=656580 $Y=779260
X4201 3333 2 3803 655 1 NR2 $T=661540 870360 0 0 $X=661540 $Y=869980
X4202 3333 2 3836 671 1 NR2 $T=669600 880440 1 0 $X=669600 $Y=875020
X4203 686 2 690 3491 1 NR2 $T=682620 779640 0 0 $X=682620 $Y=779260
X4204 3173 2 3972 655 1 NR2 $T=691920 870360 0 0 $X=691920 $Y=869980
X4205 4047 2 3902 3791 1 NR2 $T=706180 779640 0 180 $X=704320 $Y=774220
X4206 4088 2 4101 671 1 NR2 $T=713000 880440 0 180 $X=711140 $Y=875020
X4207 3234 2 4104 749 1 NR2 $T=714860 779640 1 0 $X=714860 $Y=774220
X4208 4047 2 4118 3491 1 NR2 $T=718580 789720 1 0 $X=718580 $Y=784300
X4209 3414 2 4146 749 1 NR2 $T=723540 789720 0 180 $X=721680 $Y=784300
X4210 765 2 4112 4174 1 NR2 $T=725400 729240 0 0 $X=725400 $Y=728860
X4211 766 2 4160 3498 1 NR2 $T=727260 890520 0 180 $X=725400 $Y=885100
X4212 4162 2 4155 748 1 NR2 $T=727260 749400 0 0 $X=727260 $Y=749020
X4213 3414 2 4170 748 1 NR2 $T=727260 779640 1 0 $X=727260 $Y=774220
X4214 776 2 3240 3208 1 NR2 $T=730360 789720 0 180 $X=728500 $Y=784300
X4215 774 2 777 4183 1 NR2 $T=729120 759480 0 0 $X=729120 $Y=759100
X4216 776 2 4173 4174 1 NR2 $T=732220 739320 0 180 $X=730360 $Y=733900
X4217 771 2 4182 4201 1 NR2 $T=730980 729240 0 0 $X=730980 $Y=728860
X4218 4181 2 771 4190 1 NR2 $T=732220 749400 0 0 $X=732220 $Y=749020
X4219 460 2 4148 4174 1 NR2 $T=734700 729240 0 180 $X=732840 $Y=723820
X4220 4190 2 4186 4201 1 NR2 $T=732840 749400 1 0 $X=732840 $Y=743980
X4221 4191 2 4199 774 1 NR2 $T=735940 749400 1 180 $X=734080 $Y=749020
X4222 4232 2 4218 4211 1 NR2 $T=739660 779640 0 180 $X=737800 $Y=774220
X4223 4232 2 4219 4202 1 NR2 $T=739660 799800 0 180 $X=737800 $Y=794380
X4224 4250 2 802 803 1 NR2 $T=743380 739320 0 180 $X=741520 $Y=733900
X4225 799 2 4189 4252 1 NR2 $T=741520 779640 1 0 $X=741520 $Y=774220
X4226 4255 2 4195 4211 1 NR2 $T=744000 779640 1 180 $X=742140 $Y=779260
X4227 546 2 4251 4201 1 NR2 $T=742760 749400 0 0 $X=742760 $Y=749020
X4228 4263 2 4203 4255 1 NR2 $T=745240 739320 0 180 $X=743380 $Y=733900
X4229 806 2 4196 4252 1 NR2 $T=743380 769560 0 0 $X=743380 $Y=769180
X4230 4255 2 4256 4202 1 NR2 $T=745240 789720 1 180 $X=743380 $Y=789340
X4231 3165 2 4236 4174 1 NR2 $T=744620 819960 0 0 $X=744620 $Y=819580
X4232 4255 2 4272 4209 1 NR2 $T=745240 779640 0 0 $X=745240 $Y=779260
X4233 4255 2 4267 4230 1 NR2 $T=745240 789720 1 0 $X=745240 $Y=784300
X4234 4285 2 4278 795 1 NR2 $T=750200 729240 1 180 $X=748340 $Y=728860
X4235 4280 2 4282 4230 1 NR2 $T=750200 789720 0 180 $X=748340 $Y=784300
X4236 4280 2 4288 4211 1 NR2 $T=749580 779640 1 0 $X=749580 $Y=774220
X4237 4280 2 4289 4202 1 NR2 $T=749580 789720 0 0 $X=749580 $Y=789340
X4238 4280 2 4294 4209 1 NR2 $T=750200 779640 0 0 $X=750200 $Y=779260
X4239 816 2 4292 4285 1 NR2 $T=750820 729240 0 0 $X=750820 $Y=728860
X4240 458 2 4204 828 1 NR2 $T=752060 840120 1 0 $X=752060 $Y=834700
X4241 830 2 4107 4252 1 NR2 $T=755160 769560 1 180 $X=753300 $Y=769180
X4242 4212 2 4308 4311 1 NR2 $T=753920 759480 0 0 $X=753920 $Y=759100
X4243 4315 2 4316 4211 1 NR2 $T=755780 779640 0 180 $X=753920 $Y=774220
X4244 4315 2 4303 4209 1 NR2 $T=755780 779640 1 180 $X=753920 $Y=779260
X4245 4315 2 4310 4230 1 NR2 $T=755780 789720 1 180 $X=753920 $Y=789340
X4246 4315 2 4290 4202 1 NR2 $T=755780 799800 0 180 $X=753920 $Y=794380
X4247 772 2 4322 828 1 NR2 $T=753920 840120 0 0 $X=753920 $Y=839740
X4248 812 2 4329 4315 1 NR2 $T=758880 779640 0 180 $X=757020 $Y=774220
X4249 4323 2 4324 4285 1 NR2 $T=759500 739320 0 180 $X=757640 $Y=733900
X4250 4284 2 4350 4332 1 NR2 $T=761360 769560 0 0 $X=761360 $Y=769180
X4251 4250 2 4353 840 1 NR2 $T=764460 749400 1 180 $X=762600 $Y=749020
X4252 4271 2 4372 4332 1 NR2 $T=766320 769560 1 180 $X=764460 $Y=769180
X4253 4284 2 4348 4367 1 NR2 $T=765700 769560 1 0 $X=765700 $Y=764140
X4254 4328 2 4378 4326 1 NR2 $T=767560 739320 1 0 $X=767560 $Y=733900
X4255 837 2 4379 4384 1 NR2 $T=767560 749400 0 0 $X=767560 $Y=749020
X4256 847 2 4402 4384 1 NR2 $T=768180 759480 0 0 $X=768180 $Y=759100
X4257 4328 2 4387 4386 1 NR2 $T=769420 739320 0 0 $X=769420 $Y=738940
X4258 4188 2 857 4252 1 NR2 $T=771280 789720 0 180 $X=769420 $Y=784300
X4259 4252 2 4396 3791 1 NR2 $T=770040 779640 1 0 $X=770040 $Y=774220
X4260 859 2 4399 4384 1 NR2 $T=773140 749400 1 180 $X=771280 $Y=749020
X4261 4327 2 4408 4174 1 NR2 $T=773760 769560 1 180 $X=771900 $Y=769180
X4262 772 2 4424 868 1 NR2 $T=775000 860280 1 0 $X=775000 $Y=854860
X4263 4327 2 4428 3208 1 NR2 $T=778720 789720 0 180 $X=776860 $Y=784300
X4264 458 2 4555 907 1 NR2 $T=796700 850200 0 0 $X=796700 $Y=849820
X4265 772 2 4564 907 1 NR2 $T=797940 870360 1 0 $X=797940 $Y=864940
X4266 806 2 4495 4047 1 NR2 $T=801660 779640 1 0 $X=801660 $Y=774220
X4267 830 2 4581 4047 1 NR2 $T=805380 779640 0 180 $X=803520 $Y=774220
X4268 4088 2 4605 868 1 NR2 $T=803520 870360 1 0 $X=803520 $Y=864940
X4269 4655 2 4642 929 1 NR2 $T=812200 779640 1 180 $X=810340 $Y=779260
X4270 776 2 4656 4662 1 NR2 $T=812200 749400 0 0 $X=812200 $Y=749020
X4271 4665 2 4675 4420 1 NR2 $T=815300 789720 0 0 $X=815300 $Y=789340
X4272 936 2 4680 4423 1 NR2 $T=817780 850200 0 180 $X=815920 $Y=844780
X4273 460 2 4704 4662 1 NR2 $T=817780 739320 1 0 $X=817780 $Y=733900
X4274 765 2 4738 929 1 NR2 $T=826460 789720 0 180 $X=824600 $Y=784300
X4275 4088 2 4706 828 1 NR2 $T=824600 880440 1 0 $X=824600 $Y=875020
X4276 957 2 4789 4662 1 NR2 $T=835760 739320 1 180 $X=833900 $Y=738940
X4277 4327 2 4810 4662 1 NR2 $T=840100 799800 0 180 $X=838240 $Y=794380
X4278 3165 2 4876 965 1 NR2 $T=851880 840120 1 0 $X=851880 $Y=834700
X4279 4681 2 4895 965 1 NR2 $T=852500 860280 1 0 $X=852500 $Y=854860
X4280 4657 2 4884 965 1 NR2 $T=854980 860280 1 180 $X=853120 $Y=859900
X4281 460 2 5177 5162 1 NR2 $T=904580 769560 1 0 $X=904580 $Y=764140
X4282 4655 2 5231 5162 1 NR2 $T=916980 789720 1 0 $X=916980 $Y=784300
X4283 3165 2 5244 1042 1 NR2 $T=918840 840120 0 0 $X=918840 $Y=839740
X4284 957 2 5252 5162 1 NR2 $T=923180 769560 1 180 $X=921320 $Y=769180
X4285 4327 2 5250 5162 1 NR2 $T=923180 799800 0 180 $X=921320 $Y=794380
X4286 806 2 5257 4345 1 NR2 $T=923180 769560 0 0 $X=923180 $Y=769180
X4287 4681 2 5262 1042 1 NR2 $T=925660 860280 0 180 $X=923800 $Y=854860
X4288 4088 2 5263 1042 1 NR2 $T=923800 860280 0 0 $X=923800 $Y=859900
X4289 4657 2 5331 1042 1 NR2 $T=935580 880440 1 0 $X=935580 $Y=875020
X4290 859 2 5326 4345 1 NR2 $T=942400 749400 0 0 $X=942400 $Y=749020
X4291 862 2 5309 4345 1 NR2 $T=943020 759480 0 0 $X=943020 $Y=759100
X4292 830 2 5385 4345 1 NR2 $T=943640 769560 1 0 $X=943640 $Y=764140
X4293 856 2 5649 5644 1 NR2 $T=990140 769560 0 0 $X=990140 $Y=769180
X4294 865 2 5663 5644 1 NR2 $T=995720 769560 1 180 $X=993860 $Y=769180
X4295 4681 2 5655 1113 1 NR2 $T=993860 860280 0 0 $X=993860 $Y=859900
X4296 865 2 5674 5572 1 NR2 $T=995100 779640 0 0 $X=995100 $Y=779260
X4297 5644 2 5678 963 1 NR2 $T=998820 769560 1 180 $X=996960 $Y=769180
X4298 856 2 5687 5572 1 NR2 $T=996960 779640 1 0 $X=996960 $Y=774220
X4299 5572 2 5681 963 1 NR2 $T=999440 769560 0 180 $X=997580 $Y=764140
X4300 4655 2 5691 1104 1 NR2 $T=1000060 759480 0 180 $X=998200 $Y=754060
X4301 836 2 5704 5572 1 NR2 $T=998820 739320 0 0 $X=998820 $Y=738940
X4302 836 2 5689 5644 1 NR2 $T=998820 749400 1 0 $X=998820 $Y=743980
X4303 957 2 5711 1104 1 NR2 $T=999440 769560 1 0 $X=999440 $Y=764140
X4304 4655 2 5729 892 1 NR2 $T=1001300 789720 0 0 $X=1001300 $Y=789340
X4305 4657 2 5849 1117 1 NR2 $T=1026100 890520 0 0 $X=1026100 $Y=890140
X4306 4657 2 5869 1159 1 NR2 $T=1026720 880440 0 0 $X=1026720 $Y=880060
X4307 4657 2 5891 1169 1 NR2 $T=1031060 860280 0 0 $X=1031060 $Y=859900
X4308 1922 7 1 2 INV12CK $T=326120 809880 0 0 $X=326120 $Y=809500
X4309 1922 1935 1 2 INV12CK $T=341620 819960 0 0 $X=341620 $Y=819580
X4310 2133 348 1 2 INV12CK $T=443300 860280 0 0 $X=443300 $Y=859900
X4311 348 2796 1 2 INV12CK $T=489180 860280 0 0 $X=489180 $Y=859900
X4312 3533 393 1 2 INV12CK $T=606980 759480 0 180 $X=597060 $Y=754060
X4313 3533 3314 1 2 INV12CK $T=627440 799800 0 0 $X=627440 $Y=799420
X4314 643 3533 1 2 INV12CK $T=655340 819960 0 180 $X=645420 $Y=814540
X4315 3533 622 1 2 INV12CK $T=659060 799800 0 0 $X=659060 $Y=799420
X4316 811 550 1 2 INV12CK $T=745860 729240 0 180 $X=735940 $Y=723820
X4317 811 761 1 2 INV12CK $T=785540 729240 0 180 $X=775620 $Y=723820
X4318 811 4151 1 2 INV12CK $T=785540 739320 0 180 $X=775620 $Y=733900
X4319 4631 760 1 2 INV12CK $T=808480 890520 0 180 $X=798560 $Y=885100
X4320 4631 937 1 2 INV12CK $T=822120 890520 0 0 $X=822120 $Y=890140
X4321 5312 4850 1 2 INV12CK $T=931860 840120 0 0 $X=931860 $Y=839740
X4322 5312 5317 1 2 INV12CK $T=951080 870360 0 180 $X=941160 $Y=864940
X4323 5312 1045 1 2 INV12CK $T=952320 860280 0 180 $X=942400 $Y=854860
X4324 6073 5765 1 2 INV12CK $T=1073220 850200 0 180 $X=1063300 $Y=844780
X4325 6073 1146 1 2 INV12CK $T=1070120 860280 1 0 $X=1070120 $Y=854860
X4326 1348 1307 2 1 1321 OR2 $T=230020 860280 0 180 $X=227540 $Y=854860
X4327 19 14 2 1 1376 OR2 $T=232500 739320 0 180 $X=230020 $Y=733900
X4328 24 23 2 1 1398 OR2 $T=237460 729240 0 180 $X=234980 $Y=723820
X4329 25 26 2 1 1443 OR2 $T=238700 729240 0 0 $X=238700 $Y=728860
X4330 1432 1431 2 1 1472 OR2 $T=238700 850200 1 0 $X=238700 $Y=844780
X4331 1395 1486 2 1 1498 OR2 $T=247380 819960 1 0 $X=247380 $Y=814540
X4332 1449 1520 2 1 1515 OR2 $T=254820 830040 0 180 $X=252340 $Y=824620
X4333 1567 1706 2 1 1719 OR2 $T=284580 799800 0 0 $X=284580 $Y=799420
X4334 1760 1517 2 1 1733 OR2 $T=295740 799800 1 180 $X=293260 $Y=799420
X4335 1816 1744 2 1 1802 OR2 $T=305040 789720 1 180 $X=302560 $Y=789340
X4336 1615 1854 2 1 1820 OR2 $T=313100 809880 1 180 $X=310620 $Y=809500
X4337 190 194 2 1 1843 OR2 $T=341620 880440 1 0 $X=341620 $Y=875020
X4338 2257 2227 2 1 2282 OR2 $T=375100 830040 0 0 $X=375100 $Y=829660
X4339 237 2506 2 1 2453 OR2 $T=416640 840120 1 180 $X=414160 $Y=839740
X4340 449 3165 2 1 3095 OR2 $T=537540 860280 0 180 $X=535060 $Y=854860
X4341 449 3173 2 1 437 OR2 $T=536920 880440 1 0 $X=536920 $Y=875020
X4342 452 458 2 1 3068 OR2 $T=546220 860280 0 180 $X=543740 $Y=854860
X4343 3177 460 2 1 2937 OR2 $T=548080 809880 0 180 $X=545600 $Y=804460
X4344 3177 3234 2 1 3004 OR2 $T=553660 799800 0 180 $X=551180 $Y=794380
X4345 471 3173 2 1 466 OR2 $T=554280 880440 0 0 $X=554280 $Y=880060
X4346 502 3234 2 1 3190 OR2 $T=574740 789720 0 180 $X=572260 $Y=784300
X4347 502 3414 2 1 506 OR2 $T=583420 729240 1 180 $X=580940 $Y=728860
X4348 519 3414 2 1 3252 OR2 $T=584040 739320 0 180 $X=581560 $Y=733900
X4349 520 3333 2 1 3370 OR2 $T=584040 880440 0 180 $X=581560 $Y=875020
X4350 519 3234 2 1 524 OR2 $T=584660 749400 1 0 $X=584660 $Y=743980
X4351 471 3333 2 1 3428 OR2 $T=584660 870360 1 0 $X=584660 $Y=864940
X4352 3486 3480 2 1 3301 OR2 $T=599540 789720 1 180 $X=597060 $Y=789340
X4353 4182 762 2 1 767 OR2 $T=731600 729240 0 180 $X=729120 $Y=723820
X4354 4183 4181 2 1 784 OR2 $T=731600 769560 0 0 $X=731600 $Y=769180
X4355 4181 4191 2 1 4034 OR2 $T=732220 759480 0 0 $X=732220 $Y=759100
X4356 4185 782 2 1 4202 OR2 $T=732220 789720 1 0 $X=732220 $Y=784300
X4357 782 4034 2 1 4211 OR2 $T=734080 779640 1 0 $X=734080 $Y=774220
X4358 782 784 2 1 4209 OR2 $T=734080 779640 0 0 $X=734080 $Y=779260
X4359 782 4179 2 1 4230 OR2 $T=735940 789720 0 0 $X=735940 $Y=789340
X4360 799 3480 2 1 4226 OR2 $T=742140 779640 1 180 $X=739660 $Y=779260
X4361 4232 812 2 1 3791 OR2 $T=744620 779640 1 0 $X=744620 $Y=774220
X4362 4276 4271 2 1 4232 OR2 $T=747720 769560 1 180 $X=745240 $Y=769180
X4363 4276 4284 2 1 4280 OR2 $T=750820 769560 1 180 $X=748340 $Y=769180
X4364 4300 4284 2 1 4255 OR2 $T=753300 769560 1 180 $X=750820 $Y=769180
X4365 4314 816 2 1 4242 OR2 $T=755780 739320 0 180 $X=753300 $Y=733900
X4366 4271 4300 2 1 4315 OR2 $T=755160 769560 0 0 $X=755160 $Y=769180
X4367 840 4242 2 1 835 OR2 $T=762600 739320 0 180 $X=760120 $Y=733900
X4368 816 4302 2 1 4366 OR2 $T=760120 749400 1 0 $X=760120 $Y=743980
X4369 4302 4347 2 1 842 OR2 $T=761360 729240 1 0 $X=761360 $Y=723820
X4370 4345 4334 2 1 4250 OR2 $T=761980 759480 1 0 $X=761980 $Y=754060
X4371 4302 4314 2 1 4365 OR2 $T=762600 739320 1 0 $X=762600 $Y=733900
X4372 4328 4347 2 1 4263 OR2 $T=765700 729240 1 0 $X=765700 $Y=723820
X4373 4334 4222 2 1 4367 OR2 $T=765700 759480 0 0 $X=765700 $Y=759100
X4374 843 4323 2 1 4386 OR2 $T=767560 729240 0 0 $X=767560 $Y=728860
X4375 4367 4271 2 1 4388 OR2 $T=767560 769560 1 0 $X=767560 $Y=764140
X4376 855 4263 2 1 3208 OR2 $T=768180 729240 1 0 $X=768180 $Y=723820
X4377 3791 4355 2 1 4409 OR2 $T=771280 779640 0 0 $X=771280 $Y=779260
X4378 3208 765 2 1 4391 OR2 $T=773760 789720 0 180 $X=771280 $Y=784300
X4379 835 842 2 1 519 OR2 $T=773140 729240 1 0 $X=773140 $Y=723820
X4380 841 4263 2 1 502 OR2 $T=774380 729240 0 0 $X=774380 $Y=728860
X4381 4188 4355 2 1 871 OR2 $T=774380 789720 1 0 $X=774380 $Y=784300
X4382 835 4263 2 1 475 OR2 $T=776860 729240 0 0 $X=776860 $Y=728860
X4383 841 4463 2 1 885 OR2 $T=781820 729240 0 0 $X=781820 $Y=728860
X4384 855 4463 2 1 892 OR2 $T=785540 729240 1 0 $X=785540 $Y=723820
X4385 835 4463 2 1 4312 OR2 $T=785540 739320 1 0 $X=785540 $Y=733900
X4386 965 4088 2 1 4878 OR2 $T=853740 880440 0 180 $X=851260 $Y=875020
X4387 4312 957 2 1 5671 OR2 $T=996960 799800 0 0 $X=996960 $Y=799420
X4388 885 4655 2 1 5677 OR2 $T=998820 749400 0 0 $X=998820 $Y=749020
X4389 892 957 2 1 5665 OR2 $T=998820 789720 0 0 $X=998820 $Y=789340
X4390 4312 4655 2 1 5701 OR2 $T=999440 799800 0 0 $X=999440 $Y=799420
X4391 1113 4657 2 1 5735 OR2 $T=1009360 860280 1 0 $X=1009360 $Y=854860
X4392 1117 4681 2 1 5904 OR2 $T=1030440 890520 1 0 $X=1030440 $Y=885100
X4393 1159 4681 2 1 5794 OR2 $T=1031060 880440 1 0 $X=1031060 $Y=875020
X4394 1169 4681 2 1 5923 OR2 $T=1034160 860280 1 0 $X=1034160 $Y=854860
X4395 1515 1511 1 2 1524 AN2 $T=252340 830040 0 0 $X=252340 $Y=829660
X4396 37 45 1 2 1521 AN2 $T=252960 860280 0 0 $X=252960 $Y=859900
X4397 47 1607 1 2 1646 AN2 $T=273420 890520 1 0 $X=273420 $Y=885100
X4398 1868 1893 1 2 1924 AN2 $T=326740 870360 0 0 $X=326740 $Y=869980
X4399 243 2053 1 2 2285 AN2 $T=376960 860280 0 0 $X=376960 $Y=859900
X4400 2282 2278 1 2 2307 AN2 $T=380680 830040 0 0 $X=380680 $Y=829660
X4401 4490 2 4506 4521 4018 1 NR3 $T=789260 769560 1 0 $X=789260 $Y=764140
X4402 4509 2 4525 4530 4060 1 NR3 $T=791120 769560 0 0 $X=791120 $Y=769180
X4403 4538 2 4529 4553 4022 1 NR3 $T=794220 779640 1 0 $X=794220 $Y=774220
X4404 4572 2 4587 4595 4102 1 NR3 $T=800420 860280 0 0 $X=800420 $Y=859900
X4405 921 2 4613 4618 4205 1 NR3 $T=804760 870360 0 0 $X=804760 $Y=869980
X4406 4612 2 4623 4626 4030 1 NR3 $T=806000 779640 1 0 $X=806000 $Y=774220
X4407 4516 2 4621 4630 4164 1 NR3 $T=806000 840120 0 0 $X=806000 $Y=839740
X4408 4547 2 4667 4674 4115 1 NR3 $T=813440 880440 0 0 $X=813440 $Y=880060
X4409 4602 2 4684 4689 4078 1 NR3 $T=815920 880440 1 0 $X=815920 $Y=875020
X4410 4627 2 4685 4686 4175 1 NR3 $T=815920 890520 1 0 $X=815920 $Y=885100
X4411 4756 2 4766 4790 4240 1 NR3 $T=832660 779640 1 0 $X=832660 $Y=774220
X4412 4883 2 4891 975 3991 1 NR3 $T=852500 739320 0 0 $X=852500 $Y=738940
X4413 974 2 4892 4872 4053 1 NR3 $T=852500 759480 1 0 $X=852500 $Y=754060
X4414 4931 2 4947 982 3967 1 NR3 $T=861180 759480 1 0 $X=861180 $Y=754060
X4415 5026 2 5032 1005 3913 1 NR3 $T=879780 749400 1 0 $X=879780 $Y=743980
X4416 5114 2 5122 1024 3889 1 NR3 $T=894040 749400 0 0 $X=894040 $Y=749020
X4417 1110 5686 1 5706 2 OR2B1S $T=998820 840120 1 0 $X=998820 $Y=834700
X4418 5890 5875 1 5860 2 OR2B1S $T=1031680 850200 0 180 $X=1028580 $Y=844780
X4419 3174 3074 2 1 3213 401 3099 3084 3180 453 3146 1306 ICV_7 $T=540020 749400 1 0 $X=540020 $Y=743980
X4420 3765 3662 2 1 3781 3713 3739 3735 3736 626 3723 1306 ICV_7 $T=649760 749400 0 0 $X=649760 $Y=749020
X4421 3950 3832 2 1 4028 3946 3785 3888 3965 3949 3917 1306 ICV_7 $T=693780 799800 1 0 $X=693780 $Y=794380
X4422 4001 3867 2 1 4032 3946 3898 3902 3969 3977 710 1306 ICV_7 $T=694400 779640 1 0 $X=694400 $Y=774220
X4423 739 3947 2 1 4106 4048 3898 3842 4052 4058 736 1306 ICV_7 $T=705560 769560 0 0 $X=705560 $Y=769180
X4424 4131 754 2 1 4152 728 4035 4014 3995 4124 4092 1306 ICV_7 $T=714240 880440 1 0 $X=714240 $Y=875020
X4425 4133 4009 2 1 4153 676 4035 4014 4110 4121 3821 1306 ICV_7 $T=715480 860280 1 0 $X=715480 $Y=854860
X4426 4991 4801 2 1 5005 5008 4739 4802 4964 4938 4932 1306 ICV_7 $T=868620 789720 1 0 $X=868620 $Y=784300
X4427 5093 4916 2 1 5113 5096 4915 4912 5064 5065 5053 1306 ICV_7 $T=885980 840120 1 0 $X=885980 $Y=834700
X4428 1019 4903 2 1 5107 1026 4908 4893 5088 1016 5098 1306 ICV_7 $T=889080 759480 0 0 $X=889080 $Y=759100
X4429 4997 4910 2 1 5174 5095 4982 4981 5057 4969 5136 1306 ICV_7 $T=896520 860280 0 0 $X=896520 $Y=859900
X4430 5152 964 2 1 5180 5179 4890 4918 5128 5137 5140 1306 ICV_7 $T=897140 739320 1 0 $X=897140 $Y=733900
X4431 5168 960 2 1 5192 1035 4890 4918 5145 5149 5160 1306 ICV_7 $T=899620 729240 0 0 $X=899620 $Y=728860
X4432 5447 5338 2 1 5477 1064 5326 5355 5416 5442 5405 1306 ICV_7 $T=949840 749400 0 0 $X=949840 $Y=749020
X4433 5555 5285 2 1 5584 5581 5445 5307 5526 5524 5525 1306 ICV_7 $T=967200 830040 0 0 $X=967200 $Y=829660
X4434 5596 5379 2 1 5616 5557 5328 5316 5562 5542 5583 1306 ICV_7 $T=972780 799800 1 0 $X=972780 $Y=794380
X4435 5553 5338 2 1 5625 5600 5475 5355 5577 5588 5580 1306 ICV_7 $T=974640 749400 0 0 $X=974640 $Y=749020
X4436 6221 6024 2 1 6241 6148 6147 5998 6199 6172 6207 1306 ICV_7 $T=1088720 850200 0 0 $X=1088720 $Y=849820
X4437 1232 1205 2 1 6271 6148 1227 1226 6216 1229 1228 1306 ICV_7 $T=1093680 900600 1 0 $X=1093680 $Y=895180
X4438 6338 6024 2 1 6361 6081 6147 5998 6282 6299 1245 1306 ICV_7 $T=1107940 870360 1 0 $X=1107940 $Y=864940
X4439 1248 6036 2 1 6364 1251 6109 1236 6285 6316 6324 1306 ICV_7 $T=1107940 890520 1 0 $X=1107940 $Y=885100
X4440 2499 1 2 2527 2578 1935 2164 2053 1306 ICV_8 $T=412300 830040 1 0 $X=412300 $Y=824620
X4441 2668 1 2 2705 2753 1935 2697 2565 1306 ICV_8 $T=445780 819960 0 0 $X=445780 $Y=819580
X4442 2811 1 2 2807 2838 2796 2782 2811 1306 ICV_8 $T=471200 789720 0 0 $X=471200 $Y=789340
X4443 2881 1 2 2940 2991 2796 2902 2954 1306 ICV_8 $T=494760 779640 1 0 $X=494760 $Y=774220
X4444 3146 1 2 3174 3213 393 3118 3146 1306 ICV_8 $T=533820 739320 0 0 $X=533820 $Y=738940
X4445 3455 1 2 3462 3493 3314 3510 3465 1306 ICV_8 $T=594580 840120 0 0 $X=594580 $Y=839740
X4446 3776 1 2 3801 3787 622 3750 648 1306 ICV_8 $T=656580 809880 1 0 $X=656580 $Y=804460
X4447 4068 1 2 4149 4165 760 3951 4121 1306 ICV_8 $T=717960 850200 0 0 $X=717960 $Y=849820
X4448 4103 1 2 4133 4158 760 3951 756 1306 ICV_8 $T=719820 850200 1 0 $X=719820 $Y=844780
X4449 4392 1 2 4398 4489 761 875 870 1306 ICV_8 $T=770660 749400 1 0 $X=770660 $Y=743980
X4450 4719 1 2 4751 4804 937 4712 4531 1306 ICV_8 $T=823980 870360 0 0 $X=823980 $Y=869980
X4451 4774 1 2 4803 4851 4850 4741 4805 1306 ICV_8 $T=832660 809880 0 0 $X=832660 $Y=809500
X4452 4812 1 2 4843 4873 937 4839 4719 1306 ICV_8 $T=840720 850200 0 0 $X=840720 $Y=849820
X4453 4932 1 2 4949 5001 4850 4847 4932 1306 ICV_8 $T=861180 769560 0 0 $X=861180 $Y=769180
X4454 5022 1 2 5043 5113 4850 5021 5053 1306 ICV_8 $T=878540 830040 1 0 $X=878540 $Y=824620
X4455 5087 1 2 5127 5180 4850 5034 5137 1306 ICV_8 $T=895280 749400 1 0 $X=895280 $Y=743980
X4456 5155 1 2 5205 5215 4850 5117 5203 1306 ICV_8 $T=907060 819960 0 0 $X=907060 $Y=819580
X4457 1061 1 2 5376 5450 1043 5294 5386 1306 ICV_8 $T=939300 729240 0 0 $X=939300 $Y=728860
X4458 5530 1 2 5521 5619 5317 5608 5532 1306 ICV_8 $T=974640 779640 0 0 $X=974640 $Y=779260
X4459 5931 1 2 5945 5995 1150 5974 1182 1306 ICV_8 $T=1037260 749400 1 0 $X=1037260 $Y=743980
X4460 5952 1 2 5976 5977 5765 5943 5967 1306 ICV_8 $T=1041600 840120 1 0 $X=1041600 $Y=834700
X4461 5957 1 2 5961 6005 1146 1183 5981 1306 ICV_8 $T=1042220 870360 1 0 $X=1042220 $Y=864940
X4462 5973 1 2 6012 6080 1150 5974 6032 1306 ICV_8 $T=1050900 739320 0 0 $X=1050900 $Y=738940
X4463 6103 1 2 6126 6181 5765 6140 6129 1306 ICV_8 $T=1070120 799800 1 0 $X=1070120 $Y=794380
X4464 6319 1 2 6334 6354 1150 6369 6322 1306 ICV_8 $T=1111660 749400 1 0 $X=1111660 $Y=743980
X4465 2998 2874 2 1 2994 3015 2879 2929 2969 2979 2988 1306 ICV_9 $T=502820 799800 0 0 $X=502820 $Y=799420
X4466 3098 3074 2 1 3163 428 3099 3084 3116 445 3075 1306 ICV_9 $T=531340 749400 1 0 $X=531340 $Y=743980
X4467 3426 3432 2 1 3443 3285 3404 3408 3378 3312 3399 1306 ICV_9 $T=582800 819960 1 0 $X=582800 $Y=814540
X4468 3462 3432 2 1 3488 3482 3404 3408 3450 3398 3455 1306 ICV_9 $T=591480 830040 0 0 $X=591480 $Y=829660
X4469 3474 3432 2 1 3493 3467 3401 3408 3453 3353 3465 1306 ICV_9 $T=592720 850200 1 0 $X=592720 $Y=844780
X4470 3481 538 2 1 3548 557 547 3461 3415 3423 2549 1306 ICV_9 $T=602640 880440 0 0 $X=602640 $Y=880060
X4471 3856 3832 2 1 3899 3829 3773 3748 3844 3861 3831 1306 ICV_9 $T=673320 799800 0 0 $X=673320 $Y=799420
X4472 4079 722 2 1 4105 752 4035 730 3959 4070 4072 1306 ICV_9 $T=706800 900600 1 0 $X=706800 $Y=895180
X4473 4119 3822 2 1 4134 3211 4033 661 4093 744 746 1306 ICV_9 $T=712380 739320 0 0 $X=712380 $Y=738940
X4474 4141 4127 2 1 4156 3877 4118 4014 4080 756 4103 1306 ICV_9 $T=716720 840120 0 0 $X=716720 $Y=839740
X4475 4210 4176 2 1 4239 3877 4189 4196 4138 4200 4206 1306 ICV_9 $T=732220 840120 1 0 $X=732220 $Y=834700
X4476 4215 804 2 1 4261 681 790 793 3966 796 4187 1306 ICV_9 $T=737180 890520 0 0 $X=737180 $Y=890140
X4477 4995 4801 2 1 5011 5010 4968 4802 4974 4980 4906 1306 ICV_9 $T=869860 809880 1 0 $X=869860 $Y=804460
X4478 5090 4830 2 1 5109 1020 4915 4912 5078 5047 5084 1306 ICV_9 $T=886600 870360 0 0 $X=886600 $Y=869980
X4479 5426 5393 2 1 5450 1035 5295 5287 5397 1069 5386 1306 ICV_9 $T=946120 739320 0 0 $X=946120 $Y=738940
X4480 5471 5285 2 1 5495 5195 5445 5307 5446 5432 5440 1306 ICV_9 $T=953560 830040 1 0 $X=953560 $Y=824620
X4481 5539 5393 2 1 5561 1080 5461 5287 5514 1092 5534 1306 ICV_9 $T=965340 739320 1 0 $X=965340 $Y=733900
X4482 1102 5393 2 1 5614 1074 5461 5528 5567 1099 1100 1306 ICV_9 $T=973400 739320 1 0 $X=973400 $Y=733900
X4483 6012 5803 2 1 6031 1192 5778 5946 5988 5973 1191 1306 ICV_9 $T=1049660 739320 1 0 $X=1049660 $Y=733900
X4484 6195 6153 2 1 6180 1220 5970 6178 6179 6186 6163 1306 ICV_9 $T=1085000 759480 1 0 $X=1085000 $Y=754060
X4485 6217 6104 2 1 6237 6098 6099 6136 6060 6205 6196 1306 ICV_9 $T=1088720 799800 0 0 $X=1088720 $Y=799420
X4486 6262 6104 2 1 6278 6273 6099 6136 6243 6228 6254 1306 ICV_9 $T=1096780 799800 0 0 $X=1096780 $Y=799420
X4487 6270 6091 2 1 6294 6293 6248 6178 6231 6261 6249 1306 ICV_9 $T=1098640 759480 1 0 $X=1098640 $Y=754060
X4488 6303 6026 2 1 6327 6273 6108 6100 6275 6290 6296 1306 ICV_9 $T=1103600 840120 1 0 $X=1103600 $Y=834700
X4489 6308 6104 2 1 6337 1187 6099 6136 6284 6307 6302 1306 ICV_9 $T=1104840 799800 0 0 $X=1104840 $Y=799420
X4490 6325 6093 2 1 6347 6065 6194 6069 6306 6313 6317 1306 ICV_9 $T=1107320 769560 0 0 $X=1107320 $Y=769180
X4491 6326 6084 2 1 6348 1187 6194 6069 6305 6315 6220 1306 ICV_9 $T=1107320 779640 1 0 $X=1107320 $Y=774220
X4492 2247 1 2 2513 2542 1935 2164 2247 1306 ICV_10 $T=420980 819960 1 180 $X=409200 $Y=819580
X4493 2847 1 2 2815 2813 258 2710 2778 1306 ICV_10 $T=479260 880440 0 180 $X=467480 $Y=875020
X4494 3023 1 2 3073 3080 2796 3034 3023 1306 ICV_10 $T=523280 860280 1 180 $X=511500 $Y=859900
X4495 3235 1 2 3226 3231 2796 3041 3184 1306 ICV_10 $T=552420 840120 0 180 $X=540640 $Y=834700
X4496 479 1 2 487 477 457 3141 464 1306 ICV_10 $T=559860 900600 0 180 $X=548080 $Y=895180
X4497 3612 1 2 3632 3645 3314 3644 3612 1306 ICV_10 $T=637360 789720 0 180 $X=625580 $Y=784300
X4498 4070 1 2 4137 4152 760 4123 4124 1306 ICV_10 $T=728500 870360 1 180 $X=716720 $Y=869980
X4499 4568 1 2 4615 4635 760 4583 4584 1306 ICV_10 $T=812820 860280 0 180 $X=801040 $Y=854860
X4500 4795 1 2 4816 4784 4151 4576 4726 1306 ICV_10 $T=835760 779640 1 180 $X=823980 $Y=779260
X4501 5015 1 2 5013 5007 933 4806 4952 1306 ICV_10 $T=877920 739320 1 180 $X=866140 $Y=738940
X4502 5170 1 2 5210 5207 937 5194 5157 1306 ICV_10 $T=916360 870360 0 180 $X=904580 $Y=864940
X4503 5053 1 2 5093 5425 5317 5226 5348 1306 ICV_10 $T=949840 830040 1 180 $X=938060 $Y=829660
X4504 5366 1 2 5349 5408 5317 5454 5396 1306 ICV_10 $T=963480 809880 0 180 $X=951700 $Y=804460
X4505 5432 1 2 5470 5495 5317 5337 5440 1306 ICV_10 $T=964720 819960 1 180 $X=952940 $Y=819580
X4506 5543 1 2 5586 5541 5317 5536 5482 1306 ICV_10 $T=980220 870360 1 180 $X=968440 $Y=869980
X4507 5551 1 2 5508 5616 5317 5564 5583 1306 ICV_10 $T=992000 799800 1 180 $X=980220 $Y=799420
X4508 6256 1 2 6289 6268 1146 6251 6223 1306 ICV_10 $T=1107320 860280 1 180 $X=1095540 $Y=859900
X4509 2559 1 2 2579 2585 1935 2620 2639 1306 ICV_11 $T=424080 799800 0 0 $X=424080 $Y=799420
X4510 2565 1 2 2588 2594 1935 2632 2427 1306 ICV_11 $T=425320 830040 0 0 $X=425320 $Y=829660
X4511 381 1 2 389 2864 393 392 400 1306 ICV_11 $T=477400 729240 0 0 $X=477400 $Y=728860
X4512 2899 1 2 2913 2922 2796 2966 2899 1306 ICV_11 $T=489800 840120 1 0 $X=489800 $Y=834700
X4513 2916 1 2 2925 2941 393 2986 407 1306 ICV_11 $T=492900 739320 0 0 $X=492900 $Y=738940
X4514 3051 1 2 3086 3097 2796 3141 3126 1306 ICV_11 $T=519560 850200 1 0 $X=519560 $Y=844780
X4515 3269 1 2 3344 3365 3314 3419 3364 1306 ICV_11 $T=570400 789720 0 0 $X=570400 $Y=789340
X4516 3469 1 2 3499 3505 550 3544 3469 1306 ICV_11 $T=596440 729240 0 0 $X=596440 $Y=728860
X4517 3574 1 2 3603 3604 3314 3555 3552 1306 ICV_11 $T=616280 819960 1 0 $X=616280 $Y=814540
X4518 3651 1 2 3666 3671 3314 3657 630 1306 ICV_11 $T=629300 840120 1 0 $X=629300 $Y=834700
X4519 3821 1 2 3838 3843 622 3837 3905 1306 ICV_11 $T=665260 860280 1 0 $X=665260 $Y=854860
X4520 3845 1 2 3852 3883 622 3887 3949 1306 ICV_11 $T=673320 789720 0 0 $X=673320 $Y=789340
X4521 3944 1 2 3971 4000 622 3955 4076 1306 ICV_11 $T=693160 840120 1 0 $X=693160 $Y=834700
X4522 4111 1 2 4157 4140 4151 4192 745 1306 ICV_11 $T=720440 830040 1 0 $X=720440 $Y=824620
X4523 4325 1 2 4346 4351 760 4382 4373 1306 ICV_11 $T=757020 840120 0 0 $X=757020 $Y=839740
X4524 4369 1 2 4377 4405 760 4382 882 1306 ICV_11 $T=766940 840120 1 0 $X=766940 $Y=834700
X4525 854 1 2 4414 4413 760 4461 4482 1306 ICV_11 $T=768180 880440 0 0 $X=768180 $Y=880060
X4526 4368 1 2 4403 4441 4151 4224 4456 1306 ICV_11 $T=771280 799800 1 0 $X=771280 $Y=794380
X4527 4438 1 2 4451 4534 760 4583 886 1306 ICV_11 $T=788020 840120 0 0 $X=788020 $Y=839740
X4528 5245 1 2 5284 5292 4850 5226 5366 1306 ICV_11 $T=924420 840120 1 0 $X=924420 $Y=834700
X4529 1079 1 2 5476 5487 1045 1070 1095 1306 ICV_11 $T=954800 900600 1 0 $X=954800 $Y=895180
X4530 5456 1 2 5502 5529 5317 5568 5449 1306 ICV_11 $T=962240 769560 0 0 $X=962240 $Y=769180
X4531 5588 1 2 5604 5636 1043 1109 5612 1306 ICV_11 $T=981460 739320 0 0 $X=981460 $Y=738940
X4532 1139 1 2 5807 5813 1150 5853 5841 1306 ICV_11 $T=1012460 749400 0 0 $X=1012460 $Y=749020
X4533 1154 1 2 1158 5867 5317 5819 5907 1306 ICV_11 $T=1022380 769560 0 0 $X=1022380 $Y=769180
X4534 6078 1 2 6105 6124 5765 6128 6171 1306 ICV_11 $T=1068260 840120 1 0 $X=1068260 $Y=834700
X4535 6133 1 2 6119 6158 5765 6127 6172 1306 ICV_11 $T=1075700 850200 1 0 $X=1075700 $Y=844780
X4536 2638 2 2667 1 2675 1935 2667 2598 1306 ICV_12 $T=445160 799800 0 0 $X=445160 $Y=799420
X4537 424 2 2902 1 3017 2796 3041 3037 1306 ICV_12 $T=509020 809880 0 0 $X=509020 $Y=809500
X4538 204 2 2963 1 3193 2796 3223 3182 1306 ICV_12 $T=541260 789720 1 0 $X=541260 $Y=784300
X4539 2963 2 415 1 3203 2796 3157 3235 1306 ICV_12 $T=543120 819960 1 0 $X=543120 $Y=814540
X4540 1690 2 273 1 3243 2796 3283 3264 1306 ICV_12 $T=551800 809880 1 0 $X=551800 $Y=804460
X4541 3290 2 3291 1 3340 3314 3397 3386 1306 ICV_12 $T=571020 870360 1 0 $X=571020 $Y=864940
X4542 4408 2 4422 1 4426 4151 4467 4447 1306 ICV_12 $T=773760 769560 1 0 $X=773760 $Y=764140
X4543 639 2 925 1 4620 761 934 4574 1306 ICV_12 $T=807860 729240 1 0 $X=807860 $Y=723820
X4544 4266 2 927 1 4641 760 4461 4705 1306 ICV_12 $T=807860 870360 0 0 $X=807860 $Y=869980
X4545 4738 2 4777 1 4796 4151 4576 4836 1306 ICV_12 $T=834520 789720 0 0 $X=834520 $Y=789340
X4546 4884 2 4822 1 4877 937 4927 4472 1306 ICV_12 $T=853740 870360 1 0 $X=853740 $Y=864940
X4547 973 2 5242 1 5247 4850 5226 5245 1306 ICV_12 $T=919460 830040 0 0 $X=919460 $Y=829660
X4548 5263 2 5266 1 5272 1045 5194 5350 1306 ICV_12 $T=925660 860280 0 0 $X=925660 $Y=859900
X4549 5374 2 5403 1 5404 5317 5452 5453 1306 ICV_12 $T=945500 769560 1 0 $X=945500 $Y=764140
X4550 4901 2 1085 1 5492 1045 5536 5483 1306 ICV_12 $T=959140 880440 0 0 $X=959140 $Y=880060
X4551 5691 2 5700 1 5712 5317 1135 5768 1306 ICV_12 $T=1000060 759480 1 0 $X=1000060 $Y=754060
X4552 5735 2 5782 1 5787 5317 5657 5806 1306 ICV_12 $T=1011840 850200 0 0 $X=1011840 $Y=849820
X4553 5996 2 6004 1 6029 5765 6004 6078 1306 ICV_12 $T=1053380 819960 0 0 $X=1053380 $Y=819580
X4554 6116 2 6127 1 6131 5765 6127 6165 1306 ICV_12 $T=1073840 819960 0 0 $X=1073840 $Y=819580
X4555 6168 2 6178 1 6180 5765 6224 6186 1306 ICV_12 $T=1084380 759480 0 0 $X=1084380 $Y=759100
X4556 2672 2680 2 1 2587 338 2700 2690 2688 2669 2645 1306 ICV_13 $T=446400 830040 0 180 $X=442060 $Y=824620
X4557 2745 2717 2 1 2726 2649 2756 361 2771 2716 2720 1306 ICV_13 $T=459420 870360 0 180 $X=455080 $Y=864940
X4558 2890 2874 2 1 2869 2871 2879 2739 2910 2892 2884 1306 ICV_13 $T=488560 799800 1 180 $X=484220 $Y=799420
X4559 422 2933 2 1 2941 2831 2951 2931 3022 2718 421 1306 ICV_13 $T=509020 749400 0 180 $X=504680 $Y=743980
X4560 2636 2773 2 1 2927 2871 3053 3021 3050 2610 3023 1306 ICV_13 $T=515220 850200 1 180 $X=510880 $Y=849820
X4561 3070 3074 2 1 3025 409 3099 3084 3033 3042 3076 1306 ICV_13 $T=521420 749400 0 180 $X=517080 $Y=743980
X4562 3806 3706 2 1 3774 3692 3796 3608 3833 647 3780 1306 ICV_13 $T=666500 769560 1 180 $X=662160 $Y=769180
X4563 3874 672 2 1 675 625 3896 687 3891 683 684 1306 ICV_13 $T=677040 900600 0 180 $X=672700 $Y=895180
X4564 3827 3858 2 1 3866 681 3896 3903 3907 3726 3810 1306 ICV_13 $T=679520 890520 1 180 $X=675180 $Y=890140
X4565 4109 4009 2 1 4000 3877 4118 4107 4132 4117 4076 1306 ICV_13 $T=714860 840120 0 180 $X=710520 $Y=834700
X4566 4221 4180 2 1 4172 4198 790 793 4003 4231 4214 1306 ICV_13 $T=737800 870360 0 180 $X=733460 $Y=864940
X4567 4403 4391 2 1 4319 4349 4400 4412 4419 853 4368 1306 ICV_13 $T=771900 789720 1 180 $X=767560 $Y=789340
X4568 4479 4491 2 1 4458 4357 4474 4485 4496 4478 4488 1306 ICV_13 $T=784920 850200 1 180 $X=780580 $Y=849820
X4569 4604 4575 2 1 4614 923 4427 4399 4672 4571 4597 1306 ICV_13 $T=810340 769560 0 180 $X=806000 $Y=764140
X4570 4992 4830 2 1 4951 4970 4915 4912 5012 5000 4993 1306 ICV_13 $T=873580 870360 1 180 $X=869240 $Y=869980
X4571 5043 4916 2 1 4988 5016 4915 4912 5058 4936 5022 1306 ICV_13 $T=882260 840120 0 180 $X=877920 $Y=834700
X4572 5284 5256 2 1 5247 5185 1051 5293 5296 5245 5216 1306 ICV_13 $T=928140 840120 1 180 $X=923800 $Y=839740
X4573 5278 5233 2 1 5214 1046 5295 5287 5302 5265 5255 1306 ICV_13 $T=928760 739320 1 180 $X=924420 $Y=738940
X4574 5298 5297 2 1 5219 5261 5332 5324 5335 5270 5264 1306 ICV_13 $T=931860 880440 0 180 $X=927520 $Y=875020
X4575 1065 5266 2 1 5340 5234 1067 1063 5395 1066 1068 1306 ICV_13 $T=942400 890520 1 180 $X=938060 $Y=890140
X4576 5448 5403 2 1 5413 1071 5475 5355 5480 5456 5451 1306 ICV_13 $T=954180 759480 0 180 $X=949840 $Y=754060
X4577 5552 5338 2 1 5485 5497 5475 5355 5578 5550 5449 1306 ICV_13 $T=971540 759480 0 180 $X=967200 $Y=754060
X4578 6189 6041 2 1 6166 6148 6109 6162 6202 6185 6193 1306 ICV_13 $T=1087480 880440 0 180 $X=1083140 $Y=875020
X4579 1224 1195 2 1 6159 6102 1227 1226 6187 1225 1207 1306 ICV_13 $T=1088100 890520 1 180 $X=1083760 $Y=890140
X4580 6197 6026 2 1 6124 6150 6108 6100 6209 6204 6171 1306 ICV_13 $T=1089340 840120 0 180 $X=1085000 $Y=834700
X4581 3092 1 2 3189 3132 3178 1306 ICV_14 $T=538780 870360 1 0 $X=538780 $Y=864940
X4582 3253 1 2 3318 3278 3299 1306 ICV_14 $T=559860 870360 0 0 $X=559860 $Y=869980
X4583 3118 1 2 490 3273 3275 1306 ICV_14 $T=560480 739320 1 0 $X=560480 $Y=733900
X4584 502 1 2 471 3334 3358 1306 ICV_14 $T=571020 809880 1 0 $X=571020 $Y=804460
X4585 3196 1 2 3385 3312 3339 1306 ICV_14 $T=571020 830040 0 0 $X=571020 $Y=829660
X4586 3825 1 2 672 3814 3834 1306 ICV_14 $T=663400 870360 0 0 $X=663400 $Y=869980
X4587 692 1 2 3956 3849 3830 1306 ICV_14 $T=686340 880440 0 0 $X=686340 $Y=880060
X4588 717 1 2 3946 708 716 1306 ICV_14 $T=691920 729240 1 0 $X=691920 $Y=723820
X4589 4180 1 2 804 4214 4221 1306 ICV_14 $T=736560 870360 0 0 $X=736560 $Y=869980
X4590 4435 1 2 4448 4456 4484 1306 ICV_14 $T=780580 789720 1 0 $X=780580 $Y=784300
X4591 888 1 2 923 4571 4604 1306 ICV_14 $T=798560 769560 1 0 $X=798560 $Y=764140
X4592 772 1 2 4657 4584 4610 1306 ICV_14 $T=805380 870360 1 0 $X=805380 $Y=864940
X4593 4645 1 2 4580 4637 4664 1306 ICV_14 $T=809100 729240 0 0 $X=809100 $Y=728860
X4594 4768 1 2 4778 4744 4759 1306 ICV_14 $T=833280 729240 1 0 $X=833280 $Y=723820
X4595 4814 1 2 4840 4737 4792 1306 ICV_14 $T=837620 870360 1 0 $X=837620 $Y=864940
X4596 4798 1 2 4914 971 976 1306 ICV_14 $T=850020 890520 1 0 $X=850020 $Y=885100
X4597 5257 1 2 4212 5235 5243 1306 ICV_14 $T=919460 769560 1 0 $X=919460 $Y=764140
X4598 5407 1 2 5383 5348 5392 1306 ICV_14 $T=944880 819960 1 0 $X=944880 $Y=814540
X4599 5361 1 2 5452 5449 5486 1306 ICV_14 $T=954800 769560 0 0 $X=954800 $Y=769180
X4600 5519 1 2 5541 5483 5504 1306 ICV_14 $T=962860 870360 1 0 $X=962860 $Y=864940
X4601 5454 1 2 5564 5583 5596 1306 ICV_14 $T=975880 809880 0 0 $X=975880 $Y=809500
X4602 1183 1 2 6017 6008 6040 1306 ICV_14 $T=1052140 890520 0 0 $X=1052140 $Y=890140
X4603 5888 1 2 6084 6054 6076 1306 ICV_14 $T=1060200 779640 1 0 $X=1060200 $Y=774220
X4604 5910 1 2 6093 6056 6057 1306 ICV_14 $T=1061440 789720 0 0 $X=1061440 $Y=789340
X4605 5803 1 2 1202 1196 1200 1306 ICV_14 $T=1065160 729240 1 0 $X=1065160 $Y=723820
X4606 5878 1 2 6153 6120 6142 1306 ICV_14 $T=1073840 749400 0 0 $X=1073840 $Y=749020
X4607 1394 1 2 5 1328 7 1371 8 1306 ICV_15 $T=221340 739320 0 0 $X=221340 $Y=738940
X4608 2639 1 2 2648 2590 1935 2620 2619 1306 ICV_15 $T=429660 789720 0 0 $X=429660 $Y=789340
X4609 2943 1 2 2917 2901 2796 2930 2943 1306 ICV_15 $T=488560 819960 0 0 $X=488560 $Y=819580
X4610 3009 1 2 2996 2968 393 2986 3009 1306 ICV_15 $T=502200 759480 1 0 $X=502200 $Y=754060
X4611 3048 1 2 3036 2994 2796 2947 3027 1306 ICV_15 $T=505920 799800 1 0 $X=505920 $Y=794380
X4612 3160 1 2 3159 3096 393 2986 3160 1306 ICV_15 $T=524520 759480 1 0 $X=524520 $Y=754060
X4613 464 1 2 476 455 457 3141 463 1306 ICV_15 $T=541880 890520 0 0 $X=541880 $Y=890140
X4614 3114 1 2 3123 3377 3314 3283 3334 1306 ICV_15 $T=577220 799800 0 0 $X=577220 $Y=799420
X4615 3569 1 2 3591 3539 3314 3430 2642 1306 ICV_15 $T=606980 789720 0 0 $X=606980 $Y=789340
X4616 3793 1 2 3777 3752 622 3667 3793 1306 ICV_15 $T=651620 890520 1 0 $X=651620 $Y=885100
X4617 4072 1 2 4079 4011 622 3951 3821 1306 ICV_15 $T=699360 850200 0 0 $X=699360 $Y=849820
X4618 4091 1 2 4075 4020 622 3955 4089 1306 ICV_15 $T=700600 830040 1 0 $X=700600 $Y=824620
X4619 4092 1 2 4062 4025 622 725 4092 1306 ICV_15 $T=701220 880440 0 0 $X=701220 $Y=880060
X4620 4248 1 2 4213 4177 760 3951 4248 1306 ICV_15 $T=730360 860280 0 0 $X=730360 $Y=859900
X4621 4249 1 2 4259 4287 760 822 4343 1306 ICV_15 $T=750200 880440 0 0 $X=750200 $Y=880060
X4622 4470 1 2 4460 4421 4151 4382 4470 1306 ICV_15 $T=773760 819960 0 0 $X=773760 $Y=819580
X4623 4478 1 2 4523 4458 760 4330 4488 1306 ICV_15 $T=780580 860280 1 0 $X=780580 $Y=854860
X4624 4726 1 2 4771 4679 4151 4725 4714 1306 ICV_15 $T=815920 779640 1 0 $X=815920 $Y=774220
X4625 4934 1 2 4924 4885 933 4806 4922 1306 ICV_15 $T=852500 749400 1 0 $X=852500 $Y=743980
X4626 5039 1 2 5040 4978 4850 5021 5039 1306 ICV_15 $T=870480 819960 0 0 $X=870480 $Y=819580
X4627 4938 1 2 4991 5014 4850 5042 5060 1306 ICV_15 $T=877300 779640 0 0 $X=877300 $Y=779260
X4628 5098 1 2 5071 5045 4850 4948 5098 1306 ICV_15 $T=884120 769560 1 0 $X=884120 $Y=764140
X4629 5451 1 2 5448 5413 5317 5452 5451 1306 ICV_15 $T=947360 759480 0 0 $X=947360 $Y=759100
X4630 5347 1 2 5409 5628 5317 5639 5647 1306 ICV_15 $T=982700 819960 1 0 $X=982700 $Y=814540
X4631 5645 1 2 5727 5664 1045 1107 5719 1306 ICV_15 $T=993860 870360 0 0 $X=993860 $Y=869980
X4632 5457 1 2 5490 5713 5317 5766 1127 1306 ICV_15 $T=1001300 819960 1 0 $X=1001300 $Y=814540
X4633 6164 1 2 6170 6130 5765 6088 6164 1306 ICV_15 $T=1075080 789720 1 0 $X=1075080 $Y=784300
X4634 134 2 1911 1 94 164 1306 ICV_16 $T=324880 880440 0 0 $X=324880 $Y=880060
X4635 183 2 2001 1 185 2000 1306 ICV_16 $T=336040 789720 0 0 $X=336040 $Y=789340
X4636 2053 2 2484 1 1860 2349 1306 ICV_16 $T=417880 819960 1 0 $X=417880 $Y=814540
X4637 2223 2 2171 1 2583 2545 1306 ICV_16 $T=432760 860280 1 0 $X=432760 $Y=854860
X4638 2199 2 2794 1 2199 365 1306 ICV_16 $T=467480 799800 1 0 $X=467480 $Y=794380
X4639 2930 2 3049 1 3049 3041 1306 ICV_16 $T=516460 819960 0 0 $X=516460 $Y=819580
X4640 2986 2 3128 1 3128 3118 1306 ICV_16 $T=529480 729240 0 0 $X=529480 $Y=728860
X4641 2160 2 3151 1 2160 411 1306 ICV_16 $T=533820 789720 0 0 $X=533820 $Y=789340
X4642 3233 2 3268 1 3268 474 1306 ICV_16 $T=558000 729240 1 0 $X=558000 $Y=723820
X4643 3295 2 3253 1 2949 3295 1306 ICV_16 $T=562960 870360 1 0 $X=562960 $Y=864940
X4644 3404 2 3410 1 3410 3210 1306 ICV_16 $T=580320 779640 1 0 $X=580320 $Y=774220
X4645 3485 2 3553 1 3553 3546 1306 ICV_16 $T=610700 880440 0 0 $X=610700 $Y=880060
X4646 3655 2 3680 1 3680 3669 1306 ICV_16 $T=636120 870360 0 0 $X=636120 $Y=869980
X4647 4253 2 809 1 4256 4253 1306 ICV_16 $T=742760 799800 1 0 $X=742760 $Y=794380
X4648 4316 2 4327 1 4329 4188 1306 ICV_16 $T=757020 779640 0 0 $X=757020 $Y=779260
X4649 4386 2 4389 1 4263 4395 1306 ICV_16 $T=769420 739320 1 0 $X=769420 $Y=733900
X4650 4475 2 4551 1 4551 912 1306 ICV_16 $T=797320 900600 1 0 $X=797320 $Y=895180
X4651 5326 2 5431 1 5431 5328 1306 ICV_16 $T=949840 799800 1 0 $X=949840 $Y=794380
X4652 1176 2 5876 1 1152 5941 1306 ICV_16 $T=1039120 850200 0 0 $X=1039120 $Y=849820
X4653 5564 2 5996 1 5996 6003 1306 ICV_16 $T=1048420 819960 0 0 $X=1048420 $Y=819580
X4654 5778 2 6058 1 6058 6064 1306 ICV_16 $T=1060200 739320 1 0 $X=1060200 $Y=733900
X4655 2133 1922 1 2 INV6CK $T=355260 819960 0 0 $X=355260 $Y=819580
X4656 317 2133 1 2 INV6CK $T=429660 880440 0 0 $X=429660 $Y=880060
X4657 945 4631 1 2 INV6CK $T=824600 880440 0 180 $X=819020 $Y=875020
X4658 945 6073 1 2 INV6CK $T=1065160 860280 0 180 $X=1059580 $Y=854860
X4659 3943 996 5003 5019 2 1 NR3H $T=874200 850200 0 0 $X=874200 $Y=849820
X4660 4013 998 5009 4979 2 1 NR3H $T=874820 850200 1 0 $X=874820 $Y=844780
X4661 3974 1000 5031 5033 2 1 NR3H $T=876680 840120 0 0 $X=876680 $Y=839740
X4662 3940 1004 5056 5059 2 1 NR3H $T=880400 850200 1 0 $X=880400 $Y=844780
X4663 3996 1015 5067 5055 2 1 NR3H $T=889080 880440 1 180 $X=883500 $Y=880060
X4664 3911 5176 1039 5217 2 1 NR3H $T=910160 759480 1 0 $X=910160 $Y=754060
X4665 1804 1798 1820 1 2 ND2 $T=304420 809880 0 0 $X=304420 $Y=809500
X4666 141 1865 1872 1 2 ND2 $T=316820 739320 1 0 $X=316820 $Y=733900
X4667 1986 2019 2039 1 2 ND2 $T=343480 890520 0 0 $X=343480 $Y=890140
X4668 2060 2070 2052 1 2 ND2 $T=347200 870360 1 180 $X=345340 $Y=869980
X4669 2067 2127 2114 1 2 ND2 $T=354020 799800 0 180 $X=352160 $Y=794380
X4670 2044 2118 2036 1 2 ND2 $T=354640 799800 1 180 $X=352780 $Y=799420
X4671 2067 2132 1975 1 2 ND2 $T=355880 799800 0 180 $X=354020 $Y=794380
X4672 2194 2196 2046 1 2 ND2 $T=367040 799800 1 180 $X=365180 $Y=799420
X4673 2820 1940 2833 1 2 ND2 $T=473060 739320 1 0 $X=473060 $Y=733900
X4674 4061 187 737 1 2 ND2 $T=707420 819960 1 0 $X=707420 $Y=814540
X4675 4314 4285 4328 1 2 ND2 $T=757020 729240 0 0 $X=757020 $Y=728860
X4676 4347 846 4328 1 2 ND2 $T=765700 729240 0 180 $X=763840 $Y=723820
X4677 5707 5732 5697 1 2 ND2 $T=1001300 840120 0 0 $X=1001300 $Y=839740
X4678 5858 5857 5802 1 2 ND2 $T=1025480 850200 0 0 $X=1025480 $Y=849820
X4679 4856 4826 871 4866 2 1 4874 OA112 $T=847540 789720 1 0 $X=847540 $Y=784300
X4680 945 5312 1 2 INV8CK $T=933720 860280 0 180 $X=926900 $Y=854860
X4681 4648 871 1 4659 4665 4660 2 OAI112HS $T=810960 789720 0 0 $X=810960 $Y=789340
X4682 714 177 3978 3973 1 2 ND3P $T=698120 860280 0 180 $X=693160 $Y=854860
X4683 723 171 4006 4024 1 2 ND3P $T=698120 850200 1 0 $X=698120 $Y=844780
X4684 1913 2 1987 1 2044 NR2P $T=343480 789720 1 180 $X=339760 $Y=789340
X4685 1913 2 1987 1 2067 NR2P $T=343480 789720 0 0 $X=343480 $Y=789340
X4686 847 2 4355 1 429 NR2P $T=766940 779640 0 180 $X=763220 $Y=774220
X4687 4366 2 4314 1 4225 NR2P $T=766320 749400 1 0 $X=766320 $Y=743980
X4688 427 3033 2970 2 2682 1 3044 AN4B1S $T=512740 749400 1 0 $X=512740 $Y=743980
X4689 430 3043 3026 2 2770 1 3055 AN4B1S $T=515220 759480 0 0 $X=515220 $Y=759100
X4690 434 3069 2957 2 2814 1 3087 AN4B1S $T=519560 759480 0 0 $X=519560 $Y=759100
X4691 440 3116 3022 2 2795 1 3112 AN4B1S $T=530720 749400 0 180 $X=526380 $Y=743980
X4692 451 3180 2936 2 2722 1 3192 AN4B1S $T=538780 749400 0 0 $X=538780 $Y=749020
X4693 472 3207 3228 2 2914 1 3229 AN4B1S $T=553660 759480 0 180 $X=549320 $Y=754060
X4694 2960 473 3254 2 2860 1 3257 AN4B1S $T=553660 749400 0 0 $X=553660 $Y=749020
X4695 484 3309 3272 2 2945 1 3322 AN4B1S $T=564200 769560 1 0 $X=564200 $Y=764140
X4696 498 3335 3300 2 2978 1 3326 AN4B1S $T=572880 769560 0 180 $X=568540 $Y=764140
X4697 3351 3361 3356 2 3062 1 3374 AN4B1S $T=573500 769560 1 0 $X=573500 $Y=764140
X4698 512 3372 3368 2 3108 1 3357 AN4B1S $T=579080 779640 0 180 $X=574740 $Y=774220
X4699 3412 3378 3274 2 3058 1 3363 AN4B1S $T=579700 819960 0 180 $X=575360 $Y=814540
X4700 3394 3379 3281 2 3018 1 3362 AN4B1S $T=579700 840120 0 180 $X=575360 $Y=834700
X4701 3329 3369 3373 2 2971 1 3395 AN4B1S $T=575360 860280 1 0 $X=575360 $Y=854860
X4702 3415 3406 3302 2 2781 1 3387 AN4B1S $T=582800 880440 1 180 $X=578460 $Y=880060
X4703 3434 3424 3331 2 3140 1 3422 AN4B1S $T=587760 860280 1 180 $X=583420 $Y=859900
X4704 3440 533 3341 2 2769 1 3429 AN4B1S $T=590860 900600 0 180 $X=586520 $Y=895180
X4705 3460 3450 3324 2 2985 1 3441 AN4B1S $T=595200 840120 0 180 $X=590860 $Y=834700
X4706 3468 3453 3348 2 3032 1 3457 AN4B1S $T=596440 850200 1 180 $X=592100 $Y=849820
X4707 3573 570 3326 2 3589 1 3600 AN4B1S $T=616280 769560 1 0 $X=616280 $Y=764140
X4708 3590 3594 3322 2 3599 1 3617 AN4B1S $T=618760 759480 1 0 $X=618760 $Y=754060
X4709 3625 3635 3374 2 3630 1 3643 AN4B1S $T=624960 769560 1 0 $X=624960 $Y=764140
X4710 3694 613 3357 2 3690 1 3683 AN4B1S $T=641080 779640 0 180 $X=636740 $Y=774220
X4711 4080 4071 3422 2 3920 1 4055 AN4B1S $T=711140 850200 0 180 $X=706800 $Y=844780
X4712 4097 4086 3441 2 3878 1 4063 AN4B1S $T=713620 830040 1 180 $X=709280 $Y=829660
X4713 4110 4100 3457 2 3884 1 4085 AN4B1S $T=715480 850200 0 180 $X=711140 $Y=844780
X4714 4120 4125 3363 2 3986 1 4135 AN4B1S $T=716100 809880 0 0 $X=716100 $Y=809500
X4715 4132 4138 3362 2 3957 1 4150 AN4B1S $T=719200 840120 1 0 $X=719200 $Y=834700
X4716 4208 4203 4199 2 783 1 779 AN4B1S $T=736560 739320 0 180 $X=732220 $Y=733900
X4717 1355 2 1387 1393 1351 1 1316 FA1S $T=232500 779640 1 180 $X=220720 $Y=779260
X4718 1356 2 1405 1410 1374 1 1317 FA1S $T=232500 789720 1 180 $X=220720 $Y=789340
X4719 1357 2 1385 1406 1320 1 1309 FA1S $T=232500 809880 0 180 $X=220720 $Y=804460
X4720 1358 2 1389 1379 1366 1 1307 FA1S $T=232500 830040 0 180 $X=220720 $Y=824620
X4721 1361 2 1392 1388 1378 1 1324 FA1S $T=233120 769560 0 180 $X=221340 $Y=764140
X4722 1346 2 1324 1381 1355 1 1419 FA1S $T=221340 769560 0 0 $X=221340 $Y=769180
X4723 1362 2 1344 1383 1372 1 1325 FA1S $T=233120 799800 0 180 $X=221340 $Y=794380
X4724 1347 2 1325 1357 1339 1 1395 FA1S $T=221340 809880 0 0 $X=221340 $Y=809500
X4725 1339 2 1365 1309 1358 1 1340 FA1S $T=221340 819960 1 0 $X=221340 $Y=814540
X4726 1349 2 1310 1334 12 1 16 FA1S $T=221340 870360 1 0 $X=221340 $Y=864940
X4727 1368 2 1399 1380 10 1 1313 FA1S $T=233740 890520 0 180 $X=221960 $Y=885100
X4728 1367 2 1426 1420 1401 1 1348 FA1S $T=237460 850200 0 180 $X=225680 $Y=844780
X4729 1401 2 1415 1424 1413 1 1352 FA1S $T=238080 840120 1 180 $X=226300 $Y=839740
X4730 1322 2 1467 1473 1450 1 1399 FA1S $T=244280 880440 1 180 $X=232500 $Y=880060
X4731 1351 2 1427 1466 1462 1 1404 FA1S $T=246140 809880 0 180 $X=234360 $Y=804460
X4732 1448 2 1480 1469 1463 1 22 FA1S $T=246140 870360 0 180 $X=234360 $Y=864940
X4733 1414 2 1448 1497 1461 1 1350 FA1S $T=246760 870360 1 180 $X=234980 $Y=869980
X4734 1442 2 1317 1362 1316 1 1494 FA1S $T=235600 789720 0 0 $X=235600 $Y=789340
X4735 1457 2 38 34 30 1 1403 FA1S $T=247380 900600 0 180 $X=235600 $Y=895180
X4736 1446 2 1478 1346 1428 1 1485 FA1S $T=236840 769560 0 0 $X=236840 $Y=769180
X4737 1468 2 1439 1554 1474 1 1428 FA1S $T=249240 769560 0 180 $X=237460 $Y=764140
X4738 1477 2 1501 1507 1484 1 1439 FA1S $T=251100 759480 1 180 $X=239320 $Y=759100
X4739 1470 2 1425 1458 1404 1 1486 FA1S $T=240560 809880 0 0 $X=240560 $Y=809500
X4740 1458 2 1434 1459 1464 1 1365 FA1S $T=240560 830040 1 0 $X=240560 $Y=824620
X4741 1475 2 1440 1361 1508 1 1523 FA1S $T=241180 779640 1 0 $X=241180 $Y=774220
X4742 1450 2 40 1529 1479 1 27 FA1S $T=252960 890520 0 180 $X=241180 $Y=885100
X4743 1508 2 1538 1491 1527 1 1481 FA1S $T=258540 789720 0 180 $X=246760 $Y=784300
X4744 1514 2 1542 1470 1494 1 1525 FA1S $T=248000 809880 1 0 $X=248000 $Y=804460
X4745 1517 2 1552 1468 1446 1 1567 FA1S $T=249240 769560 0 0 $X=249240 $Y=769180
X4746 1474 2 1356 1481 1555 1 1553 FA1S $T=249240 789720 0 0 $X=249240 $Y=789340
X4747 1518 2 1553 1442 1419 1 1563 FA1S $T=249240 799800 1 0 $X=249240 $Y=794380
X4748 1533 2 1561 1503 1543 1 1497 FA1S $T=261020 870360 1 180 $X=249240 $Y=869980
X4749 1531 2 1506 1513 1526 1 1572 FA1S $T=251720 749400 1 0 $X=251720 $Y=743980
X4750 1552 2 1597 1586 1523 1 1478 FA1S $T=264740 779640 0 180 $X=252960 $Y=774220
X4751 1586 2 1603 1617 1601 1 1381 FA1S $T=269700 779640 1 180 $X=257920 $Y=779260
X4752 1589 2 1516 1611 1602 1 1554 FA1S $T=270320 769560 0 180 $X=258540 $Y=764140
X4753 6375 2 1569 1618 1531 1 1628 FA1S $T=261020 739320 1 0 $X=261020 $Y=733900
X4754 1592 2 1566 1575 1477 1 1620 FA1S $T=261020 749400 0 0 $X=261020 $Y=749020
X4755 1308 2 1623 1647 1627 1 1583 FA1S $T=275280 870360 1 180 $X=263500 $Y=869980
X4756 1609 2 1589 1634 1620 1 1643 FA1S $T=264120 769560 0 0 $X=264120 $Y=769180
X4757 1555 2 1582 1590 1621 1 1542 FA1S $T=264120 799800 1 0 $X=264120 $Y=794380
X4758 1585 2 1660 1583 1632 1 1380 FA1S $T=279620 880440 1 180 $X=267840 $Y=880060
X4759 77 2 1663 1681 83 1 64 FA1S $T=279620 900600 0 180 $X=267840 $Y=895180
X4760 1618 2 1605 1614 1639 1 1668 FA1S $T=269080 739320 0 0 $X=269080 $Y=738940
X4761 1642 2 1572 1668 1609 1 1688 FA1S $T=270940 749400 1 0 $X=270940 $Y=743980
X4762 1634 2 1689 1633 1669 1 1597 FA1S $T=283340 779640 0 180 $X=271560 $Y=774220
X4763 1600 2 1694 1670 1676 1 73 FA1S $T=283960 890520 1 180 $X=272180 $Y=890140
X4764 1649 2 1629 1637 1656 1 1705 FA1S $T=272800 759480 0 0 $X=272800 $Y=759100
X4765 1671 2 1705 1643 1713 1 1706 FA1S $T=276520 779640 0 0 $X=276520 $Y=779260
X4766 1672 2 1680 1737 1725 1 1660 FA1S $T=291400 880440 1 180 $X=279620 $Y=880060
X4767 1702 2 1664 1684 1691 1 1741 FA1S $T=280240 769560 1 0 $X=280240 $Y=764140
X4768 6376 2 1700 1683 1665 1 1775 FA1S $T=280860 749400 0 0 $X=280860 $Y=749020
X4769 1543 2 1743 1749 1686 1 1480 FA1S $T=292640 870360 1 180 $X=280860 $Y=869980
X4770 1694 2 1697 103 1729 1 1681 FA1S $T=293260 900600 0 180 $X=281480 $Y=895180
X4771 6377 2 1673 1710 1766 1 1774 FA1S $T=285200 739320 1 0 $X=285200 $Y=733900
X4772 1731 2 1649 1702 1768 1 1716 FA1S $T=285820 759480 0 0 $X=285820 $Y=759100
X4773 1438 2 1771 1761 1759 1 1473 FA1S $T=297600 880440 0 180 $X=285820 $Y=875020
X4774 1744 2 1755 1671 1790 1 1760 FA1S $T=288300 789720 0 0 $X=288300 $Y=789340
X4775 1768 2 1778 1736 1779 1 1727 FA1S $T=301320 779640 1 180 $X=289540 $Y=779260
X4776 1755 2 1727 1741 1475 1 1713 FA1S $T=290160 789720 1 0 $X=290160 $Y=784300
X4777 6378 2 1801 1775 1818 1 1767 FA1S $T=308140 749400 1 180 $X=296360 $Y=749020
X4778 6379 2 1767 1822 1642 1 1846 FA1S $T=296980 749400 1 0 $X=296980 $Y=743980
X4779 1417 2 1817 1835 1783 1 1461 FA1S $T=309380 870360 1 180 $X=297600 $Y=869980
X4780 1430 2 124 1836 1806 1 1783 FA1S $T=309380 890520 0 180 $X=297600 $Y=885100
X4781 1815 2 1841 1850 1592 1 1722 FA1S $T=310000 769560 0 180 $X=298220 $Y=764140
X4782 1801 2 1784 1776 1808 1 1841 FA1S $T=298220 769560 0 0 $X=298220 $Y=769180
X4783 1817 2 1845 1838 1679 1 1463 FA1S $T=310000 870360 0 180 $X=298220 $Y=864940
X4784 6380 2 1774 1810 1628 1 1822 FA1S $T=299460 739320 1 0 $X=299460 $Y=733900
X4785 6381 2 1827 1731 1815 1 1853 FA1S $T=299460 759480 0 0 $X=299460 $Y=759100
X4786 1561 2 1840 125 1839 1 115 FA1S $T=311240 880440 1 180 $X=299460 $Y=880060
X4787 6382 2 1879 1875 1819 1 1810 FA1S $T=316200 789720 0 180 $X=304420 $Y=784300
X4788 1858 2 126 1864 1866 1 6383 FA1S $T=317440 789720 1 180 $X=305660 $Y=789340
X4789 1818 2 1889 1842 1887 1 1850 FA1S $T=322400 769560 1 180 $X=310620 $Y=769180
X4790 6384 2 1853 1732 1846 1 1816 FA1S $T=311240 759480 0 0 $X=311240 $Y=759100
X4791 6385 2 1874 1910 1903 1 1827 FA1S $T=325500 769560 0 180 $X=313720 $Y=764140
X4792 1675 2 1924 1914 1904 1 1835 FA1S $T=326740 870360 1 180 $X=314960 $Y=869980
X4793 1960 2 1995 2011 1974 1 1745 FA1S $T=336040 779640 0 180 $X=324260 $Y=774220
X4794 1963 2 2005 1962 1983 1 1918 FA1S $T=337280 759480 0 180 $X=325500 $Y=754060
X4795 178 2 2016 189 181 1 1928 FA1S $T=338520 729240 0 180 $X=326740 $Y=723820
X4796 1977 2 2068 1999 1960 1 1723 FA1S $T=338520 769560 1 180 $X=326740 $Y=769180
X4797 179 2 2032 1928 1992 1 1933 FA1S $T=339140 729240 1 180 $X=327360 $Y=728860
X4798 1992 2 2012 1957 1963 1 1937 FA1S $T=340380 749400 0 180 $X=328600 $Y=743980
X4799 1983 2 2057 2013 1977 1 1938 FA1S $T=340380 759480 1 180 $X=328600 $Y=759100
X4800 2012 2 2051 2033 2021 1 1962 FA1S $T=343480 749400 1 180 $X=331700 $Y=749020
X4801 2032 2 2079 2097 2028 1 1957 FA1S $T=346580 739320 0 180 $X=334800 $Y=733900
X4802 1974 2 2075 2080 2042 1 1770 FA1S $T=346580 779640 1 180 $X=334800 $Y=779260
X4803 2049 2 2088 2076 2064 1 2011 FA1S $T=349680 779640 0 180 $X=337900 $Y=774220
X4804 2055 2 2074 2087 1894 1 2010 FA1S $T=349680 890520 0 180 $X=337900 $Y=885100
X4805 2057 2 2092 2029 2049 1 1999 FA1S $T=350300 769560 0 180 $X=338520 $Y=764140
X4806 2005 2 2103 2102 2048 1 2013 FA1S $T=350920 759480 0 180 $X=339140 $Y=754060
X4807 2016 2 206 2083 2089 1 2028 FA1S $T=352160 729240 0 180 $X=340380 $Y=723820
X4808 2083 2 2128 2101 2091 1 2033 FA1S $T=353400 729240 1 180 $X=341620 $Y=728860
X4809 2066 2 2096 2010 195 1 208 FA1S $T=342240 900600 1 0 $X=342240 $Y=895180
X4810 2079 2 2124 2131 2108 1 2021 FA1S $T=354640 739320 1 180 $X=342860 $Y=738940
X4811 2006 2 2056 197 2146 1 6386 FA1S $T=344720 809880 1 0 $X=344720 $Y=804460
X4812 2051 2 2116 2159 2120 1 2048 FA1S $T=357120 749400 1 180 $X=345340 $Y=749020
X4813 2140 2 2163 2175 2018 1 201 FA1S $T=360840 890520 1 180 $X=349060 $Y=890140
X4814 2080 2 2094 2024 2154 1 1811 FA1S $T=349680 789720 1 0 $X=349680 $Y=784300
X4815 2139 2 1950 2162 2071 1 2175 FA1S $T=351540 890520 1 0 $X=351540 $Y=885100
X4816 2043 2 2122 187 2169 1 2093 FA1S $T=363940 809880 1 180 $X=352160 $Y=809500
X4817 2103 2 2176 2129 2172 1 2068 FA1S $T=364560 769560 0 180 $X=352780 $Y=764140
X4818 216 2 2178 221 2130 1 2089 FA1S $T=365800 729240 0 180 $X=354020 $Y=723820
X4819 2131 2 2192 2137 2173 1 2102 FA1S $T=365800 759480 0 180 $X=354020 $Y=754060
X4820 2064 2 2202 2145 2180 1 2042 FA1S $T=367040 779640 0 180 $X=355260 $Y=774220
X4821 220 2 2198 2205 2166 1 210 FA1S $T=367660 900600 0 180 $X=355880 $Y=895180
X4822 2146 2 2157 225 2188 1 6387 FA1S $T=368280 809880 0 180 $X=356500 $Y=804460
X4823 230 2 2179 2216 2213 1 2097 FA1S $T=372620 739320 0 180 $X=360840 $Y=733900
X4824 2216 2 2239 2249 2221 1 2108 FA1S $T=374480 749400 0 180 $X=362700 $Y=743980
X4825 234 2 2220 2224 2225 1 219 FA1S $T=374480 880440 0 180 $X=362700 $Y=875020
X4826 2220 2 2258 2261 2143 1 223 FA1S $T=375720 880440 1 180 $X=363940 $Y=880060
X4827 2173 2 2259 2237 2233 1 2029 FA1S $T=376340 749400 1 180 $X=364560 $Y=749020
X4828 2172 2 2201 2193 2231 1 1995 FA1S $T=367040 769560 1 0 $X=367040 $Y=764140
X4829 2268 2 2285 2230 2279 1 2224 FA1S $T=382540 870360 1 180 $X=370760 $Y=869980
X4830 248 2 2286 2269 2284 1 2213 FA1S $T=383160 729240 1 180 $X=371380 $Y=728860
X4831 2271 2 2241 2272 2274 1 2163 FA1S $T=373860 890520 0 0 $X=373860 $Y=890140
X4832 2280 2 2335 2266 2308 1 1943 FA1S $T=386880 779640 0 180 $X=375100 $Y=774220
X4833 2221 2 2294 2347 2333 1 2159 FA1S $T=389980 749400 0 180 $X=378200 $Y=743980
X4834 2326 2 2341 2358 2280 1 1980 FA1S $T=390600 769560 1 180 $X=378820 $Y=769180
X4835 2308 2 2359 2283 2339 1 1958 FA1S $T=390600 779640 1 180 $X=378820 $Y=779260
X4836 2335 2 2357 2363 2353 1 2283 FA1S $T=392460 759480 1 180 $X=380680 $Y=759100
X4837 2341 2 2368 2362 2298 1 2266 FA1S $T=393080 759480 0 180 $X=381300 $Y=754060
X4838 2304 2 262 2270 2313 1 2225 FA1S $T=382540 880440 1 0 $X=382540 $Y=875020
X4839 2339 2 2387 2379 2365 1 1949 FA1S $T=395560 789720 1 180 $X=383780 $Y=789340
X4840 2365 2 2336 2394 2371 1 2165 FA1S $T=396180 799800 0 180 $X=384400 $Y=794380
X4841 2284 2 2345 2338 260 1 2101 FA1S $T=387500 729240 0 0 $X=387500 $Y=728860
X4842 2359 2 2410 2366 2375 1 2379 FA1S $T=390600 779640 0 0 $X=390600 $Y=779260
X4843 2389 2 2426 2449 2417 1 2366 FA1S $T=403620 769560 1 180 $X=391840 $Y=769180
X4844 2410 2 2432 2443 2415 1 2336 FA1S $T=404240 789720 0 180 $X=392460 $Y=784300
X4845 2401 2 2428 2454 2414 1 2374 FA1S $T=404860 759480 0 180 $X=393080 $Y=754060
X4846 2357 2 2455 2380 2424 1 2375 FA1S $T=404860 769560 0 180 $X=393080 $Y=764140
X4847 2414 2 2448 2435 2407 1 2380 FA1S $T=405480 749400 0 180 $X=393700 $Y=743980
X4848 2368 2 2450 2389 2374 1 2353 FA1S $T=405480 759480 1 180 $X=393700 $Y=759100
X4849 2431 2 2472 2401 2422 1 2362 FA1S $T=407960 739320 1 180 $X=396180 $Y=738940
X4850 2387 2 2457 2463 2452 1 2394 FA1S $T=408580 789720 1 180 $X=396800 $Y=789340
X4851 2452 2 2485 2464 2460 1 2405 FA1S $T=409820 799800 1 180 $X=398040 $Y=799420
X4852 2371 2 2490 2405 2469 1 2295 FA1S $T=411060 809880 0 180 $X=399280 $Y=804460
X4853 2469 2 2480 2491 2475 1 2296 FA1S $T=412300 809880 1 180 $X=400520 $Y=809500
X4854 2288 2 2458 2026 2446 1 2500 FA1S $T=401140 880440 0 0 $X=401140 $Y=880060
X4855 2473 2 2495 2508 2481 1 2422 FA1S $T=413540 739320 0 180 $X=401760 $Y=733900
X4856 2458 2 2265 2437 2254 1 2507 FA1S $T=402380 890520 0 0 $X=402380 $Y=890140
X4857 2510 2 2462 2445 2479 1 302 FA1S $T=409820 900600 1 0 $X=409820 $Y=895180
X4858 2460 2 2504 2505 2536 1 2475 FA1S $T=412300 799800 0 0 $X=412300 $Y=799420
X4859 2417 2 2501 2518 2482 1 2463 FA1S $T=412920 769560 1 0 $X=412920 $Y=764140
X4860 2491 2 2498 2497 2517 1 2148 FA1S $T=413540 809880 1 0 $X=413540 $Y=804460
X4861 2548 2 2566 2560 2557 1 2363 FA1S $T=426560 759480 1 180 $X=414780 $Y=759100
X4862 2540 2 2529 2507 300 1 309 FA1S $T=414780 890520 1 0 $X=414780 $Y=885100
X4863 2481 2 2538 2488 303 1 2560 FA1S $T=415400 739320 1 0 $X=415400 $Y=733900
X4864 2415 2 2535 2541 2516 1 2490 FA1S $T=417880 789720 1 0 $X=417880 $Y=784300
X4865 313 2 2563 2553 310 1 2609 FA1S $T=423460 729240 0 0 $X=423460 $Y=728860
X4866 2584 2 306 2510 315 1 325 FA1S $T=424700 900600 1 0 $X=424700 $Y=895180
X4867 2595 2 2576 2431 2634 1 2612 FA1S $T=426560 749400 0 0 $X=426560 $Y=749020
X4868 2607 2 2556 328 2575 1 2576 FA1S $T=438960 739320 1 180 $X=427180 $Y=738940
X4869 2596 2 2577 316 2569 1 2635 FA1S $T=427800 759480 1 0 $X=427800 $Y=754060
X4870 2605 2 2568 2473 2609 1 2634 FA1S $T=429040 739320 1 0 $X=429040 $Y=733900
X4871 2614 2 2616 2637 2326 1 1971 FA1S $T=440820 779640 0 180 $X=429040 $Y=774220
X4872 2537 2 2584 2500 2540 1 332 FA1S $T=429040 890520 1 0 $X=429040 $Y=885100
X4873 2616 2 2626 2631 2612 1 2358 FA1S $T=441440 769560 1 180 $X=429660 $Y=769180
X4874 2626 2 2647 2548 2635 1 2298 FA1S $T=442680 759480 1 180 $X=430900 $Y=759100
X4875 2624 2 2544 323 330 1 2658 FA1S $T=433380 729240 1 0 $X=433380 $Y=723820
X4876 2659 2 2658 2673 2605 1 2625 FA1S $T=449500 729240 1 180 $X=437720 $Y=728860
X4877 2665 2 2595 2625 2653 1 2637 FA1S $T=441440 759480 1 0 $X=441440 $Y=754060
X4878 2702 2 346 2703 2713 1 2653 FA1S $T=455080 749400 0 180 $X=443300 $Y=743980
X4879 2703 2 2646 2596 2714 1 2631 FA1S $T=455080 749400 1 180 $X=443300 $Y=749020
X4880 2686 2 2663 2607 2654 1 2713 FA1S $T=443920 739320 0 0 $X=443920 $Y=738940
X4881 2715 2 2665 2728 2614 1 2030 FA1S $T=458180 769560 0 180 $X=446400 $Y=764140
X4882 354 2 351 2624 2711 1 2742 FA1S $T=448880 729240 1 0 $X=448880 $Y=723820
X4883 2758 2 2764 2763 2715 1 2599 FA1S $T=467480 759480 0 180 $X=455700 $Y=754060
X4884 2764 2 2702 2808 2779 1 2728 FA1S $T=468720 749400 0 180 $X=456940 $Y=743980
X4885 6388 2 2798 369 2758 1 2589 FA1S $T=468720 749400 1 180 $X=456940 $Y=749020
X4886 2762 2 2742 2659 372 1 2779 FA1S $T=458800 739320 1 0 $X=458800 $Y=733900
X4887 367 2 362 364 2686 1 2808 FA1S $T=460660 729240 0 0 $X=460660 $Y=728860
X4888 2798 2 2762 375 374 1 2763 FA1S $T=474920 739320 1 180 $X=463140 $Y=738940
X4889 1311 1329 1338 2 1 XNR2HS $T=220720 860280 0 0 $X=220720 $Y=859900
X4890 1345 1337 1360 2 1 XNR2HS $T=224440 880440 0 0 $X=224440 $Y=880060
X4891 1391 1386 13 2 1 XNR2HS $T=233120 870360 1 180 $X=227540 $Y=869980
X4892 1332 1430 1345 2 1 XNR2HS $T=239320 890520 0 180 $X=233740 $Y=885100
X4893 1482 1489 1502 2 1 XNR2HS $T=247380 840120 0 0 $X=247380 $Y=839740
X4894 1359 1509 1551 2 1 XNR2HS $T=254820 819960 0 0 $X=254820 $Y=819580
X4895 1648 1645 1391 2 1 XNR2HS $T=277760 870360 0 180 $X=272180 $Y=864940
X4896 1630 1666 1674 2 1 XNR2HS $T=279000 809880 1 0 $X=279000 $Y=804460
X4897 1707 1726 1746 2 1 XNR2HS $T=289540 819960 1 0 $X=289540 $Y=814540
X4898 141 1900 1902 2 1 XNR2HS $T=321160 739320 1 0 $X=321160 $Y=733900
X4899 2027 2041 2052 2 1 XNR2HS $T=341000 860280 0 0 $X=341000 $Y=859900
X4900 2222 2232 2215 2 1 XNR2HS $T=373860 809880 1 180 $X=368280 $Y=809500
X4901 2388 2323 2381 2 1 XNR2HS $T=394940 819960 1 0 $X=394940 $Y=814540
X4902 2440 2434 2386 2 1 XNR2HS $T=404860 840120 0 180 $X=399280 $Y=834700
X4903 2461 2429 2391 2 1 XNR2HS $T=405480 860280 1 0 $X=405480 $Y=854860
X4904 2537 2066 2547 2 1 XNR2HS $T=417880 890520 0 0 $X=417880 $Y=890140
X4905 2547 307 2392 2 1 XNR2HS $T=424080 890520 0 0 $X=424080 $Y=890140
X4906 4276 4250 4275 2 1 XNR2HS $T=753300 759480 0 180 $X=747720 $Y=754060
X4907 1546 1521 1510 1 2 1455 OA12 $T=256060 870360 0 180 $X=252340 $Y=864940
X4908 52 1505 1492 1 2 1496 OA12 $T=256060 880440 1 180 $X=252340 $Y=880060
X4909 1535 1591 1587 1 2 1467 OA12 $T=267220 870360 0 180 $X=263500 $Y=864940
X4910 1619 1711 1720 1 2 1734 OA12 $T=285200 809880 1 0 $X=285200 $Y=804460
X4911 2045 2112 2107 1 2 2096 OA12 $T=354020 880440 1 180 $X=350300 $Y=880060
X4912 4186 775 767 1 2 4147 OA12 $T=731600 749400 0 180 $X=727880 $Y=743980
X4913 4278 818 4268 1 2 4207 OA12 $T=749580 739320 0 180 $X=745860 $Y=733900
X4914 4276 4250 4299 1 2 4311 OA12 $T=758260 759480 0 180 $X=754540 $Y=754060
X4915 1535 1 1545 1535 1529 1558 2 OAI22S $T=256060 890520 1 0 $X=256060 $Y=885100
X4916 1860 1 1968 1965 1967 60 2 OAI22S $T=335420 870360 0 180 $X=331700 $Y=864940
X4917 2001 1 1982 1990 1934 180 2 OAI22S $T=337900 799800 0 180 $X=334180 $Y=794380
X4918 1994 1 2014 1994 2026 2017 2 OAI22S $T=337900 880440 1 0 $X=337900 $Y=875020
X4919 2820 1 379 2839 382 377 2 OAI22S $T=476780 729240 1 0 $X=476780 $Y=723820
X4920 546 4270 768 1 2 4268 AO12 $T=749580 739320 1 180 $X=745860 $Y=738940
X4921 1311 1321 2 1330 1 1318 AOI12HS $T=220100 850200 0 0 $X=220100 $Y=849820
X4922 1482 1472 2 1454 1 1377 AOI12HS $T=247380 840120 1 180 $X=243040 $Y=839740
X4923 1498 1359 2 1519 1 1536 AOI12HS $T=252960 819960 1 0 $X=252960 $Y=814540
X4924 1593 1606 2 1584 1 1619 AOI12HS $T=270320 809880 1 180 $X=265980 $Y=809500
X4925 1724 1733 2 1739 1 1720 AOI12HS $T=288920 799800 0 0 $X=288920 $Y=799420
X4926 1719 1726 2 1724 1 1754 AOI12HS $T=289540 809880 0 0 $X=289540 $Y=809500
X4927 2262 2273 2 2238 1 2276 AOI12HS $T=381300 809880 0 180 $X=376960 $Y=804460
X4928 2302 2323 2 2273 1 2264 AOI12HS $T=387500 809880 1 180 $X=383160 $Y=809500
X4929 2385 2323 2 2360 1 2364 AOI12HS $T=394320 809880 1 180 $X=389980 $Y=809500
X4930 2409 2399 2 2421 1 2303 AOI12HS $T=398660 840120 0 0 $X=398660 $Y=839740
X4931 2453 2440 2 2470 1 2372 AOI12HS $T=404860 840120 1 0 $X=404860 $Y=834700
X4932 1540 2 1594 1624 1 AN2B1S $T=269700 860280 0 0 $X=269700 $Y=859900
X4933 1662 2 1659 1591 1 AN2B1S $T=280240 860280 1 180 $X=277140 $Y=859900
X4934 1750 2 1821 1825 1 AN2B1S $T=305040 890520 0 0 $X=305040 $Y=890140
X4935 173 2 1951 1966 1 AN2B1S $T=331080 900600 1 0 $X=331080 $Y=895180
X4936 2117 2 2142 2112 1 AN2B1S $T=358360 870360 1 180 $X=355260 $Y=869980
X4937 2406 2 2412 2471 1 AN2B1S $T=404860 880440 1 0 $X=404860 $Y=875020
X4938 1318 1336 1 1353 2 1359 OAI12HS $T=224440 830040 0 0 $X=224440 $Y=829660
X4939 1377 1364 1 1354 2 1311 OAI12HS $T=230640 860280 1 180 $X=226920 $Y=859900
X4940 1530 1536 1 1550 2 1593 OAI12HS $T=262260 809880 0 0 $X=262260 $Y=809500
X4941 1570 1576 1 1571 2 1584 OAI12HS $T=266600 799800 1 180 $X=262880 $Y=799420
X4942 1565 1625 1 1570 2 1666 OAI12HS $T=275280 809880 0 0 $X=275280 $Y=809500
X4943 97 1902 1 1909 2 1917 OAI12HS $T=321780 749400 0 0 $X=321780 $Y=749020
X4944 2039 1986 1 2019 2 2027 OAI12HS $T=342240 890520 1 180 $X=338520 $Y=890140
X4945 2052 2060 1 2070 2 2078 OAI12HS $T=347200 870360 0 0 $X=347200 $Y=869980
X4946 187 2067 1 2132 2 2149 OAI12HS $T=359600 799800 0 180 $X=355880 $Y=794380
X4947 226 2194 1 2127 2 2203 OAI12HS $T=369520 789720 1 180 $X=365800 $Y=789340
X4948 157 2044 1 2196 2 2214 OAI12HS $T=371380 799800 0 180 $X=367660 $Y=794380
X4949 2243 2204 1 2210 2 2238 OAI12HS $T=375100 809880 0 180 $X=371380 $Y=804460
X4950 2263 2264 1 2243 2 2232 OAI12HS $T=378820 809880 1 180 $X=375100 $Y=809500
X4951 253 2194 1 2118 2 2277 OAI12HS $T=381920 799800 1 180 $X=378200 $Y=799420
X4952 2303 2290 1 2276 2 2169 OAI12HS $T=383160 809880 1 180 $X=379440 $Y=809500
X4953 2337 2322 1 2312 2 2273 OAI12HS $T=387500 809880 0 180 $X=383780 $Y=804460
X4954 2372 2367 1 2354 2 2399 OAI12HS $T=399280 840120 0 180 $X=395560 $Y=834700
X4955 2418 2425 1 2436 2 2421 OAI12HS $T=401140 850200 1 0 $X=401140 $Y=844780
X4956 2404 2430 1 2418 2 2429 OAI12HS $T=404860 860280 0 180 $X=401140 $Y=854860
X4957 2278 2444 1 2433 2 2440 OAI12HS $T=403000 830040 1 0 $X=403000 $Y=824620
X4958 4212 4191 1 4190 2 4229 OAI12HS $T=741520 759480 0 180 $X=737800 $Y=754060
X4959 2086 2078 1 2086 200 2078 2 MOAI1 $T=352160 880440 0 180 $X=347820 $Y=875020
X4960 2392 271 1 2392 2039 271 2 MOAI1 $T=399280 900600 0 180 $X=394940 $Y=895180
X4961 2299 1 2 2831 2807 2656 2838 2831 1306 ICV_19 $T=471200 789720 1 0 $X=471200 $Y=784300
X4962 3041 1 2 3196 3162 2965 3188 3101 1306 ICV_19 $T=537540 830040 0 0 $X=537540 $Y=829660
X4963 488 1 2 3330 3294 3287 3232 3317 1306 ICV_19 $T=562960 850200 0 0 $X=562960 $Y=849820
X4964 3875 1 2 695 688 685 696 695 1306 ICV_19 $T=679520 729240 1 0 $X=679520 $Y=723820
X4965 929 1 2 907 4615 4596 4634 4357 1306 ICV_19 $T=806000 850200 0 0 $X=806000 $Y=849820
X4966 3211 1 2 952 943 4580 949 923 1306 ICV_19 $T=822120 729240 1 0 $X=822120 $Y=723820
X4967 4385 1 2 4976 4695 4916 4962 4976 1306 ICV_19 $T=866760 840120 1 0 $X=866760 $Y=834700
X4968 5132 1 2 5189 5173 4910 5199 5096 1306 ICV_19 $T=904580 850200 1 0 $X=904580 $Y=844780
X4969 5256 1 2 5434 5392 5256 5425 4976 1306 ICV_19 $T=944880 840120 1 0 $X=944880 $Y=834700
X4970 5591 1 2 5535 5535 5304 5585 5557 1306 ICV_19 $T=972160 860280 0 0 $X=972160 $Y=859900
X4971 4976 1 2 5956 5940 5797 5912 5956 1306 ICV_19 $T=1038500 819960 0 0 $X=1038500 $Y=819580
X4972 5920 1 2 5993 5961 5926 5985 1185 1306 ICV_19 $T=1042840 860280 0 0 $X=1042840 $Y=859900
X4973 5984 1 2 6039 5997 5923 6027 1185 1306 ICV_19 $T=1050280 850200 0 0 $X=1050280 $Y=849820
X4974 1192 1 2 6018 6022 5878 6049 1192 1306 ICV_19 $T=1054620 759480 1 0 $X=1054620 $Y=754060
X4975 6067 1 2 6095 6063 5878 6080 1080 1306 ICV_19 $T=1062680 749400 0 0 $X=1062680 $Y=749020
X4976 1195 1 2 1208 6096 1145 6106 6047 1306 ICV_19 $T=1068880 890520 0 0 $X=1068880 $Y=890140
X4977 1799 7 1824 2 1 102 1738 1793 1306 ICV_20 $T=298220 830040 0 0 $X=298220 $Y=829660
X4978 2332 258 2373 2 1 2330 2310 2319 1306 ICV_20 $T=383160 860280 0 0 $X=383160 $Y=859900
X4979 3396 3314 3419 2 1 3438 3375 3389 1306 ICV_20 $T=576600 769560 0 0 $X=576600 $Y=769180
X4980 3653 3314 3687 2 1 621 3638 3646 1306 ICV_20 $T=626820 860280 0 0 $X=626820 $Y=859900
X4981 4444 760 4461 2 1 4453 4425 4432 1306 ICV_20 $T=774380 880440 1 0 $X=774380 $Y=875020
X4982 4663 760 4712 2 1 946 4649 4658 1306 ICV_20 $T=810960 860280 0 0 $X=810960 $Y=859900
X4983 5076 4850 5117 2 1 5121 5061 5068 1306 ICV_20 $T=884120 830040 0 0 $X=884120 $Y=829660
X4984 5182 937 5227 2 1 5136 5189 5186 1306 ICV_20 $T=906440 850200 0 0 $X=906440 $Y=849820
X4985 5623 1045 1108 2 1 5660 5602 5618 1306 ICV_20 $T=978980 890520 0 0 $X=978980 $Y=890140
X4986 5574 1043 1109 2 1 5606 5559 5498 1306 ICV_20 $T=981460 729240 1 0 $X=981460 $Y=723820
X4987 5769 5765 5805 2 1 5784 5754 5762 1306 ICV_20 $T=1006260 789720 1 0 $X=1006260 $Y=784300
X4988 5814 5317 5856 2 1 5844 5798 5801 1306 ICV_20 $T=1014940 819960 0 0 $X=1014940 $Y=819580
X4989 5894 1150 5853 2 1 5944 5877 5886 1306 ICV_20 $T=1029200 729240 0 0 $X=1029200 $Y=728860
X4990 5906 5765 5564 2 1 5925 5889 5898 1306 ICV_20 $T=1030440 830040 0 0 $X=1030440 $Y=829660
X4991 5947 5765 5943 2 1 5952 5835 5827 1306 ICV_20 $T=1037880 819960 1 0 $X=1037880 $Y=814540
X4992 5978 1146 6017 2 1 6016 5965 5971 1306 ICV_20 $T=1042840 890520 1 0 $X=1042840 $Y=885100
X4993 5887 1 1168 2 BUF6CK $T=1036020 739320 1 0 $X=1036020 $Y=733900
X4994 1712 2 1652 1 1781 1721 1708 1764 1717 1306 ICV_21 $T=293260 830040 0 0 $X=293260 $Y=829660
X4995 109 2 1752 1 1792 1785 1792 1785 1701 1306 ICV_21 $T=297600 860280 0 0 $X=297600 $Y=859900
X4996 1984 2 2099 1 2050 1828 2058 2115 2109 1306 ICV_21 $T=350300 830040 1 0 $X=350300 $Y=824620
X4997 2329 2 2061 1 304 2530 2522 252 2309 1306 ICV_21 $T=417260 860280 0 0 $X=417260 $Y=859900
X4998 2852 2 384 1 2684 2478 2684 384 2834 1306 ICV_21 $T=479880 870360 1 0 $X=479880 $Y=864940
X4999 2203 2 3015 1 3004 3036 3004 3003 3016 1306 ICV_21 $T=510880 799800 0 0 $X=510880 $Y=799420
X5000 3264 2 3286 1 3035 3269 3301 3286 3296 1306 ICV_21 $T=561720 799800 1 0 $X=561720 $Y=794380
X5001 3569 2 3621 1 3623 3574 582 3621 3596 1306 ICV_21 $T=622480 809880 0 0 $X=622480 $Y=809500
X5002 3691 2 3664 1 3647 620 3647 3664 3677 1306 ICV_21 $T=637980 830040 1 0 $X=637980 $Y=824620
X5003 4201 2 4270 1 4222 768 4201 4275 817 1306 ICV_21 $T=745860 749400 0 0 $X=745860 $Y=749020
X5004 768 2 4293 1 4270 4308 4293 4299 4279 1306 ICV_21 $T=750820 749400 1 0 $X=750820 $Y=743980
X5005 4390 2 4410 1 4412 4401 4409 4410 4420 1306 ICV_21 $T=772520 819960 1 0 $X=772520 $Y=814540
X5006 4373 2 4418 1 4394 4438 4409 4418 4423 1306 ICV_21 $T=773140 850200 1 0 $X=773140 $Y=844780
X5007 4428 2 4435 1 4435 876 4448 4434 4442 1306 ICV_21 $T=775620 779640 0 0 $X=775620 $Y=779260
X5008 4439 2 874 1 874 4414 874 878 4445 1306 ICV_21 $T=777480 890520 0 0 $X=777480 $Y=890140
X5009 883 2 4475 1 887 4466 887 878 4471 1306 ICV_21 $T=783060 890520 0 0 $X=783060 $Y=890140
X5010 4551 2 4556 1 903 911 903 848 4561 1306 ICV_21 $T=795460 890520 0 0 $X=795460 $Y=890140
X5011 5868 2 1162 1 5830 1171 1162 1168 1164 1306 ICV_21 $T=1029820 729240 1 0 $X=1029820 $Y=723820
X5012 5881 2 5910 1 5910 5934 5910 5887 5918 1306 ICV_21 $T=1033540 799800 1 0 $X=1033540 $Y=794380
X5013 3989 5108 1022 5077 2 1 NR3HT $T=888460 850200 1 0 $X=888460 $Y=844780
X5014 3897 5175 5211 1040 2 1 NR3HT $T=905820 749400 0 0 $X=905820 $Y=749020
X5015 4225 963 1 2 INV4CK $T=838240 759480 1 0 $X=838240 $Y=754060
X5016 834 4389 4395 2 1 4431 AN3 $T=771900 739320 1 0 $X=771900 $Y=733900
X5017 849 4323 4355 1 2 OR2P $T=765700 739320 0 0 $X=765700 $Y=738940
X5018 4365 4323 867 1 2 OR2P $T=771280 739320 0 0 $X=771280 $Y=738940
X5019 4309 836 1 2 INV3 $T=758260 739320 0 0 $X=758260 $Y=738940
X5020 4350 830 1 2 INV3 $T=760740 779640 1 0 $X=760740 $Y=774220
X5021 843 4314 1 2 INV3 $T=763840 739320 1 180 $X=761360 $Y=738940
X5022 858 856 1 2 INV3 $T=770660 729240 1 0 $X=770660 $Y=723820
X5023 4380 1 2 859 INV3CK $T=770040 759480 1 0 $X=770040 $Y=754060
X5024 1373 2 1447 1433 1 1373 1459 1396 1306 ICV_22 $T=239940 819960 0 0 $X=239940 $Y=819580
X5025 1400 2 1516 1418 1 20 1507 1532 1306 ICV_22 $T=252960 759480 1 0 $X=252960 $Y=754060
X5026 1644 2 1631 1650 1 1581 1651 1650 1306 ICV_22 $T=275900 789720 0 0 $X=275900 $Y=789340
X5027 110 2 1842 1638 1 110 1848 1704 1306 ICV_22 $T=308140 779640 1 0 $X=308140 $Y=774220
X5028 143 2 1875 1638 1 29 1874 1885 1306 ICV_22 $T=314960 779640 0 0 $X=314960 $Y=779260
X5029 2017 2 2045 184 1 151 196 1777 1306 ICV_22 $T=342860 880440 0 0 $X=342860 $Y=880060
X5030 193 2 2071 1911 1 1777 2087 203 1306 ICV_22 $T=346580 880440 0 0 $X=346580 $Y=880060
X5031 2113 2 2091 207 1 205 2120 207 1306 ICV_22 $T=352160 739320 1 0 $X=352160 $Y=733900
X5032 2084 2 2076 211 1 2113 2129 211 1306 ICV_22 $T=355260 769560 0 0 $X=355260 $Y=769180
X5033 2255 2 2269 211 1 2255 2294 2125 1306 ICV_22 $T=377580 739320 0 0 $X=377580 $Y=738940
X5034 270 2 2437 259 1 188 2462 252 1306 ICV_22 $T=403620 900600 1 0 $X=403620 $Y=895180
X5035 292 2 2450 294 1 2468 2472 294 1306 ICV_22 $T=410440 759480 1 0 $X=410440 $Y=754060
X5036 288 2 2508 286 1 287 2502 2489 1306 ICV_22 $T=412920 729240 0 0 $X=412920 $Y=728860
X5037 295 2 2538 2474 1 295 2553 286 1306 ICV_22 $T=417880 729240 0 0 $X=417880 $Y=728860
X5038 288 2 2525 293 1 301 2575 296 1306 ICV_22 $T=421600 749400 1 0 $X=421600 $Y=743980
X5039 4232 2 4241 4230 1 4232 4246 4209 1306 ICV_22 $T=739660 789720 1 0 $X=739660 $Y=784300
X5040 3480 2 4295 839 1 837 2895 4355 1306 ICV_22 $T=759500 779640 0 0 $X=759500 $Y=779260
X5041 4194 761 755 812 1 2 QDFFRBP $T=733460 739320 0 0 $X=733460 $Y=738940
X5042 820 4151 4129 4222 1 2 QDFFRBP $T=749580 759480 1 180 $X=737180 $Y=759100
X5043 4279 4151 4224 4284 1 2 QDFFRBP $T=748340 769560 1 0 $X=748340 $Y=764140
X5044 3714 4243 1 2 BUF2CK $T=740900 840120 0 0 $X=740900 $Y=839740
X5045 3870 3087 3889 3894 1 2 3890 AO13S $T=677660 759480 1 0 $X=677660 $Y=754060
X5046 3880 3112 3897 3894 1 2 3912 AO13S $T=678900 749400 0 0 $X=678900 $Y=749020
X5047 3904 3055 3911 3894 1 2 3928 AO13S $T=681380 759480 0 0 $X=681380 $Y=759100
X5048 3769 3192 3913 3894 1 2 3930 AO13S $T=682000 759480 1 0 $X=682000 $Y=754060
X5049 3933 701 3940 3941 1 2 3934 AO13S $T=686340 870360 0 0 $X=686340 $Y=869980
X5050 3942 3429 3943 3941 1 2 3916 AO13S $T=691300 890520 0 180 $X=686960 $Y=885100
X5051 3960 3044 3967 3894 1 2 3978 AO13S $T=691300 749400 0 0 $X=691300 $Y=749020
X5052 715 713 3974 3941 1 2 3871 AO13S $T=696260 890520 0 180 $X=691920 $Y=885100
X5053 3982 3257 3991 3894 1 2 4006 AO13S $T=695640 759480 1 0 $X=695640 $Y=754060
X5054 724 721 3996 3941 1 2 3973 AO13S $T=700600 890520 0 180 $X=696260 $Y=885100
X5055 4002 3395 4013 3941 1 2 4024 AO13S $T=698740 860280 1 0 $X=698740 $Y=854860
X5056 4160 4205 786 4179 1 2 4220 AO13S $T=733460 799800 0 0 $X=733460 $Y=799420
X5057 3629 4240 798 4034 1 2 4233 AO13S $T=738420 769560 0 0 $X=738420 $Y=769180
X5058 3998 726 2 541 1 ND2F $T=698740 809880 1 0 $X=698740 $Y=804460
X5059 3979 3387 3989 3941 1 2 3983 AO13 $T=695020 870360 0 0 $X=695020 $Y=869980
X5060 3912 3983 3998 1 2 AN2T $T=694400 809880 1 0 $X=694400 $Y=804460
X5061 3871 1 3890 691 2 218 ND3HT $T=675800 850200 1 0 $X=675800 $Y=844780
X5062 3916 1 3930 702 2 495 ND3HT $T=682620 819960 1 0 $X=682620 $Y=814540
X5063 3934 1 3928 707 2 237 ND3HT $T=685720 850200 0 0 $X=685720 $Y=849820
X5064 3791 686 2 1 3697 OR2S $T=679520 779640 1 180 $X=677040 $Y=779260
X5065 669 1 3846 174 2 ND2P $T=670220 819960 1 0 $X=670220 $Y=814540
X5066 670 1 3847 157 2 ND2P $T=670220 819960 0 0 $X=670220 $Y=819580
X5067 678 1 3872 3448 2 ND2P $T=674560 809880 0 0 $X=674560 $Y=809500
X5068 680 1 3873 226 2 ND2P $T=674560 819960 1 0 $X=674560 $Y=814540
X5069 311 2554 1 1940 2542 2523 2 MOAI1H $T=427800 819960 0 180 $X=420360 $Y=814540
X5070 1429 1447 1420 1 2 1397 HA1 $T=242420 850200 1 180 $X=234360 $Y=849820
X5071 1453 1422 1462 1 2 1320 HA1 $T=238080 819960 1 0 $X=238080 $Y=814540
X5072 1452 1476 1374 1 2 1372 HA1 $T=247380 799800 0 180 $X=239320 $Y=794380
X5073 35 1445 1413 1 2 1432 HA1 $T=249240 840120 0 180 $X=241180 $Y=834700
X5074 37 1488 1464 1 2 1366 HA1 $T=251100 830040 1 180 $X=243040 $Y=829660
X5075 1612 1631 1602 1 2 1601 HA1 $T=274040 789720 0 180 $X=265980 $Y=784300
X5076 1635 1651 1527 1 2 1621 HA1 $T=278380 799800 1 180 $X=270320 $Y=799420
X5077 1712 1730 1691 1 2 1669 HA1 $T=291400 769560 1 180 $X=283340 $Y=769180
X5078 1823 1848 1808 1 2 1779 HA1 $T=311240 779640 1 180 $X=303180 $Y=779260
X5079 1814 1859 6389 1 2 1819 HA1 $T=314340 799800 1 180 $X=306280 $Y=799420
X5080 1794 1862 1903 1 2 1887 HA1 $T=329840 779640 1 180 $X=321780 $Y=779260
X5081 2040 2062 2024 1 2 1781 HA1 $T=347200 789720 0 180 $X=339140 $Y=784300
X5082 2167 2187 2145 1 2 2154 HA1 $T=367040 779640 1 180 $X=358980 $Y=779260
X5083 2207 2228 2193 1 2 2180 HA1 $T=373240 769560 1 180 $X=365180 $Y=769180
X5084 2256 2267 2237 1 2 2231 HA1 $T=380060 759480 1 180 $X=372000 $Y=759100
X5085 2331 2297 2347 1 2 2233 HA1 $T=383160 749400 0 0 $X=383160 $Y=749020
X5086 2361 2346 2338 1 2 2333 HA1 $T=395560 739320 1 180 $X=387500 $Y=738940
X5087 2486 2466 2497 1 2 6390 HA1 $T=406100 779640 0 0 $X=406100 $Y=779260
X5088 2502 2524 2488 1 2 2407 HA1 $T=417880 739320 1 180 $X=409820 $Y=738940
X5089 2503 2525 2435 1 2 2482 HA1 $T=417880 749400 0 180 $X=409820 $Y=743980
X5090 2539 2526 2518 1 2 2516 HA1 $T=424080 779640 0 180 $X=416020 $Y=774220
X5091 2531 2511 2505 1 2 2517 HA1 $T=424080 799800 0 180 $X=416020 $Y=794380
X5092 2534 2564 2541 1 2 2536 HA1 $T=426560 779640 1 180 $X=418500 $Y=779260
X5093 1318 1326 1333 2 1 XOR2HS $T=220100 840120 0 0 $X=220100 $Y=839740
X5094 1377 1416 1437 2 1 XOR2HS $T=235600 860280 0 0 $X=235600 $Y=859900
X5095 1536 1539 1598 2 1 XOR2HS $T=262260 819960 1 0 $X=262260 $Y=814540
X5096 1625 1640 1657 2 1 XOR2HS $T=274660 819960 1 0 $X=274660 $Y=814540
X5097 1763 1754 1787 2 1 XOR2HS $T=295120 809880 0 0 $X=295120 $Y=809500
X5098 1780 1734 1795 2 1 XOR2HS $T=296980 799800 0 0 $X=296980 $Y=799420
X5099 2291 2264 2324 2 1 XOR2HS $T=381920 819960 1 0 $X=381920 $Y=814540
X5100 2351 2364 2340 2 1 XOR2HS $T=393080 819960 0 180 $X=387500 $Y=814540
X5101 2372 2369 2350 2 1 XOR2HS $T=393700 840120 1 180 $X=388120 $Y=839740
X5102 2278 2416 2378 2 1 XOR2HS $T=402380 830040 0 180 $X=396800 $Y=824620
X5103 2419 2430 2356 2 1 XOR2HS $T=401760 860280 0 0 $X=401760 $Y=859900
X5104 185 2194 2 171 1 2299 MUX2S $T=376340 789720 0 0 $X=376340 $Y=789340
X5105 222 2044 237 2242 1 2 MUX2P $T=370140 789720 0 0 $X=370140 $Y=789340
X5106 1722 1716 1688 1 2 1732 MAO222 $T=285200 759480 1 0 $X=285200 $Y=754060
X5107 150 143 142 1 2 1872 MAO222 $T=314960 729240 1 0 $X=314960 $Y=723820
X5108 1892 152 1897 1 2 1866 MAO222 $T=321780 799800 0 180 $X=316820 $Y=794380
X5109 1826 156 1858 1 2 1916 MAO222 $T=320540 789720 0 0 $X=320540 $Y=789340
X5110 162 160 1934 1 2 1897 MAO222 $T=327980 799800 0 180 $X=323020 $Y=794380
X5111 1917 166 1916 1 2 1981 MAO222 $T=326120 789720 0 0 $X=326120 $Y=789340
X5112 186 2000 2006 1 2 1982 MAO222 $T=339140 799800 1 180 $X=334180 $Y=799420
X5113 232 2217 2181 1 2 2188 MAO222 $T=367040 799800 0 0 $X=367040 $Y=799420
X5114 1722 1716 1688 2 1 1790 XOR3 $T=291400 759480 1 0 $X=291400 $Y=754060
X5115 131 137 155 2 1 1892 XOR3 $T=312480 779640 1 0 $X=312480 $Y=774220
X5116 174 1984 2043 2 1 2050 XOR3 $T=333560 809880 1 0 $X=333560 $Y=804460
X5117 1864 81 2 118 130 1 1788 FA1 $T=313720 729240 0 180 $X=298220 $Y=723820
X5118 1826 148 2 1888 1788 1 1900 FA1 $T=306900 729240 0 0 $X=306900 $Y=728860
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=15 FDC=0
X0 1 2 3 4 5 6 MUX2 $T=0 0 0 0 $X=0 $Y=-380
X1 7 8 9 10 4 11 3 AOI22S $T=0 0 1 180 $X=-3720 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 BUF1S $T=0 0 0 0 $X=0 $Y=-380
X1 5 6 3 2 7 8 MUX2 $T=6820 0 1 180 $X=2480 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=0
X0 1 2 3 4 5 6 MUX2 $T=-4340 0 0 0 $X=-4340 $Y=-380
X1 7 8 3 4 9 10 MUX2 $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT BUF3 I VCC GND O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN3S I1 I2 I3 GND VCC O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR3B2 I1 B1 VCC O B2 GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF4CK I GND O VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI13HS B3 O B2 B1 VCC A1 GND
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22HT A2 A1 VCC B1 O B2 GND
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MAO222P A1 B1 C1 O GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=0
X0 1 2 3 4 DELA $T=0 0 0 0 $X=0 $Y=-380
X1 5 2 3 6 DELA $T=4960 0 0 0 $X=4960 $Y=-380
.ENDS
***************************************
.SUBCKT ND2T I2 GND I1 O VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF6 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXL2HS B S OB A VCC GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HA1P A B C S GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6 7 8 9 10 11 12 13
** N=13 EP=13 IP=16 FDC=0
X0 1 2 3 4 5 6 7 OAI22S $T=0 0 0 0 $X=0 $Y=-380
X1 8 2 9 10 11 12 7 OAI22S $T=4340 0 0 0 $X=4340 $Y=-380
.ENDS
***************************************
.SUBCKT XNR3 I2 I1 I3 VCC GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540
+ 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560
+ 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580
+ 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640
+ 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660
+ 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680
+ 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700
+ 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720
+ 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740
+ 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760
+ 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780
+ 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800
+ 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820
+ 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840
+ 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860
+ 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880
+ 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900
+ 901 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920
+ 921 922 923 924 925 926 927 928 929 930 931 932 933 934 935 936 937 938 939 940
+ 941 942 943 944 945 946 947 948 949 950 951 952 953 954 955 956 957 958 959 960
+ 961 962 963 964 965 966 967 968 969 970 971 972 973 974 975 976 977 978 979 980
+ 981 982 983 984 985 986 987 988 989 990 991 992 993 994 995 996 997 998 999 1000
+ 1001 1002 1003 1004 1005 1006 1007 1008 1009 1010 1011 1012 1013 1014 1015 1016 1017 1018 1019 1020
+ 1021 1022 1023 1024 1025 1026 1027 1028 1029 1030 1031 1032 1033 1034 1035 1036 1037 1038 1039 1040
+ 1041 1042 1043 1044 1045 1046 1047 1048 1049 1050 1051 1052 1053 1054 1055 1056 1057 1058 1059 1060
+ 1061 1062 1063 1064 1065 1066 1067 1068 1069 1070 1071 1072 1073 1074 1075 1076 1077 1078 1079 1080
+ 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 1093 1094 1095 1096 1097 1098 1099 1100
+ 1101 1102 1103 1104 1105 1106 1107 1108 1109 1110 1111 1112 1113 1114 1115 1116 1117 1118 1119 1120
+ 1121 1122 1123 1124 1125 1126 1127 1128 1129 1130 1131 1132 1133 1134 1135 1136 1137 1138 1139 1140
+ 1141 1142 1143 1144 1145 1146 1147 1148 1149 1150 1151 1152 1153 1154 1155 1156 1157 1158 1159 1160
+ 1161 1162 1163 1164 1165 1166 1167 1168 1169 1170 1171 1172 1173 1174 1175 1176 1177 1178 1179 1180
+ 1181 1182 1183 1184 1185 1186 1187 1188 1189 1190 1191 1192 1193 1194 1204 1233
** N=6244 EP=1196 IP=32847 FDC=0
X0 1192 1193 1193 1193 1204 1193 1194 YA2GSD $T=1349740 530520 0 90 $X=1210240 $Y=533370
X1 3 2 1265 1 INV1S $T=220720 588120 0 0 $X=220720 $Y=587740
X2 9 2 1240 1 INV1S $T=221960 628440 0 180 $X=220720 $Y=623020
X3 1247 2 1235 1 INV1S $T=221960 638520 1 180 $X=220720 $Y=638140
X4 14 2 1263 1 INV1S $T=224440 547800 1 180 $X=223200 $Y=547420
X5 15 2 1270 1 INV1S $T=225060 648600 0 180 $X=223820 $Y=643180
X6 5 2 1254 1 INV1S $T=226920 567960 0 0 $X=226920 $Y=567580
X7 20 2 1280 1 INV1S $T=229400 658680 1 180 $X=228160 $Y=658300
X8 22 2 1287 1 INV1S $T=230020 678840 1 180 $X=228780 $Y=678460
X9 1310 2 23 1 INV1S $T=231880 719160 0 0 $X=231880 $Y=718780
X10 1272 2 1247 1 INV1S $T=233740 678840 1 0 $X=233740 $Y=673420
X11 1290 2 1321 1 INV1S $T=233740 709080 0 0 $X=233740 $Y=708700
X12 8 2 1329 1 INV1S $T=236840 598200 1 180 $X=235600 $Y=597820
X13 6 2 1327 1 INV1S $T=238080 557880 0 180 $X=236840 $Y=552460
X14 4 2 1276 1 INV1S $T=238080 608280 0 180 $X=236840 $Y=602860
X15 1350 2 1324 1 INV1S $T=240560 699000 1 180 $X=239320 $Y=698620
X16 1403 2 32 1 INV1S $T=249240 618360 1 180 $X=248000 $Y=617980
X17 1247 2 1418 1 INV1S $T=249860 638520 0 0 $X=249860 $Y=638140
X18 1387 2 1413 1 INV1S $T=254820 547800 1 180 $X=253580 $Y=547420
X19 1387 2 45 1 INV1S $T=255440 537720 1 180 $X=254200 $Y=537340
X20 41 2 1462 1 INV1S $T=256060 537720 0 0 $X=256060 $Y=537340
X21 1449 2 1430 1 INV1S $T=256060 719160 0 0 $X=256060 $Y=718780
X22 1409 2 1415 1 INV1S $T=257920 719160 0 180 $X=256680 $Y=713740
X23 1403 2 1376 1 INV1S $T=259780 567960 0 180 $X=258540 $Y=562540
X24 1408 2 1386 1 INV1S $T=258540 588120 1 0 $X=258540 $Y=582700
X25 44 2 1444 1 INV1S $T=263500 557880 0 180 $X=262260 $Y=552460
X26 49 2 1443 1 INV1S $T=263500 608280 1 180 $X=262260 $Y=607900
X27 57 2 1456 1 INV1S $T=263500 699000 0 180 $X=262260 $Y=693580
X28 1497 2 1403 1 INV1S $T=265360 588120 0 180 $X=264120 $Y=582700
X29 57 2 1501 1 INV1S $T=264740 688920 0 0 $X=264740 $Y=688540
X30 1496 2 57 1 INV1S $T=265980 699000 1 180 $X=264740 $Y=698620
X31 1485 2 1496 1 INV1S $T=269080 699000 1 180 $X=267840 $Y=698620
X32 1513 2 1539 1 INV1S $T=269080 557880 0 0 $X=269080 $Y=557500
X33 1524 2 1460 1 INV1S $T=270940 699000 1 180 $X=269700 $Y=698620
X34 66 2 68 1 INV1S $T=269700 719160 1 0 $X=269700 $Y=713740
X35 1520 2 62 1 INV1S $T=271560 547800 1 180 $X=270320 $Y=547420
X36 58 2 1514 1 INV1S $T=271560 638520 1 180 $X=270320 $Y=638140
X37 1491 2 1533 1 INV1S $T=271560 638520 0 0 $X=271560 $Y=638140
X38 1528 2 1507 1 INV1S $T=272800 567960 0 0 $X=272800 $Y=567580
X39 1539 2 74 1 INV1S $T=274040 547800 0 0 $X=274040 $Y=547420
X40 73 2 1548 1 INV1S $T=274040 578040 0 0 $X=274040 $Y=577660
X41 1552 2 1511 1 INV1S $T=276520 547800 1 180 $X=275280 $Y=547420
X42 1545 2 1556 1 INV1S $T=275280 699000 0 0 $X=275280 $Y=698620
X43 1539 2 1540 1 INV1S $T=279000 557880 0 0 $X=279000 $Y=557500
X44 1507 2 76 1 INV1S $T=280240 567960 0 180 $X=279000 $Y=562540
X45 1564 2 1571 1 INV1S $T=279620 588120 1 0 $X=279620 $Y=582700
X46 46 2 1582 1 INV1S $T=280240 578040 1 0 $X=280240 $Y=572620
X47 1571 2 73 1 INV1S $T=281480 578040 1 180 $X=280240 $Y=577660
X48 1462 2 1579 1 INV1S $T=281480 557880 1 0 $X=281480 $Y=552460
X49 1558 2 1497 1 INV1S $T=281480 588120 0 0 $X=281480 $Y=587740
X50 1578 2 1584 1 INV1S $T=282720 618360 0 180 $X=281480 $Y=612940
X51 1462 2 1604 1 INV1S $T=283340 557880 1 0 $X=283340 $Y=552460
X52 81 2 1428 1 INV1S $T=283340 699000 0 0 $X=283340 $Y=698620
X53 1509 2 1591 1 INV1S $T=286440 638520 0 180 $X=285200 $Y=633100
X54 1571 2 1616 1 INV1S $T=287060 578040 0 0 $X=287060 $Y=577660
X55 1580 2 1617 1 INV1S $T=288920 598200 0 180 $X=287680 $Y=592780
X56 1507 2 1631 1 INV1S $T=290160 567960 1 0 $X=290160 $Y=562540
X57 75 2 90 1 INV1S $T=290160 719160 1 0 $X=290160 $Y=713740
X58 80 2 91 1 INV1S $T=290780 578040 1 0 $X=290780 $Y=572620
X59 97 2 1500 1 INV1S $T=293260 709080 1 180 $X=292020 $Y=708700
X60 1454 2 97 1 INV1S $T=292640 688920 1 0 $X=292640 $Y=683500
X61 1641 2 1606 1 INV1S $T=295120 598200 0 180 $X=293880 $Y=592780
X62 1556 2 1634 1 INV1S $T=295120 688920 1 180 $X=293880 $Y=688540
X63 56 2 1454 1 INV1S $T=294500 658680 0 0 $X=294500 $Y=658300
X64 1659 2 89 1 INV1S $T=296360 567960 0 180 $X=295120 $Y=562540
X65 1661 2 94 1 INV1S $T=296360 688920 0 180 $X=295120 $Y=683500
X66 103 2 102 1 INV1S $T=297600 688920 0 180 $X=296360 $Y=683500
X67 1661 2 1464 1 INV1S $T=300080 688920 0 180 $X=298840 $Y=683500
X68 1675 2 1645 1 INV1S $T=301320 557880 1 180 $X=300080 $Y=557500
X69 1687 2 1530 1 INV1S $T=301940 578040 1 180 $X=300700 $Y=577660
X70 1634 2 55 1 INV1S $T=301940 688920 0 180 $X=300700 $Y=683500
X71 1635 2 1711 1 INV1S $T=301320 688920 0 0 $X=301320 $Y=688540
X72 1547 2 1651 1 INV1S $T=304420 668760 1 180 $X=303180 $Y=668380
X73 1657 2 109 1 INV1S $T=303180 709080 0 0 $X=303180 $Y=708700
X74 1697 2 110 1 INV1S $T=306280 719160 0 180 $X=305040 $Y=713740
X75 1654 2 1716 1 INV1S $T=306280 699000 1 0 $X=306280 $Y=693580
X76 1539 2 1720 1 INV1S $T=306900 567960 0 0 $X=306900 $Y=567580
X77 1687 2 1623 1 INV1S $T=306900 578040 0 0 $X=306900 $Y=577660
X78 1706 2 1718 1 INV1S $T=308760 688920 0 180 $X=307520 $Y=683500
X79 121 2 1687 1 INV1S $T=311240 578040 0 180 $X=310000 $Y=572620
X80 1681 2 1721 1 INV1S $T=311240 638520 1 180 $X=310000 $Y=638140
X81 117 2 118 1 INV1S $T=310000 688920 1 0 $X=310000 $Y=683500
X82 1757 2 1761 1 INV1S $T=314340 567960 1 0 $X=314340 $Y=562540
X83 1730 2 1759 1 INV1S $T=315580 588120 1 180 $X=314340 $Y=587740
X84 1766 2 1771 1 INV1S $T=315580 598200 1 0 $X=315580 $Y=592780
X85 125 2 1739 1 INV1S $T=316200 638520 0 0 $X=316200 $Y=638140
X86 1741 2 1787 1 INV1S $T=317440 598200 0 0 $X=317440 $Y=597820
X87 1786 2 1743 1 INV1S $T=319920 567960 0 180 $X=318680 $Y=562540
X88 101 2 1797 1 INV1S $T=320540 719160 0 0 $X=320540 $Y=718780
X89 1797 2 1755 1 INV1S $T=321160 688920 1 0 $X=321160 $Y=683500
X90 1805 2 1775 1 INV1S $T=323020 668760 0 180 $X=321780 $Y=663340
X91 1805 2 1809 1 INV1S $T=323020 668760 1 0 $X=323020 $Y=663340
X92 1755 2 1805 1 INV1S $T=323020 668760 0 0 $X=323020 $Y=668380
X93 1810 2 1806 1 INV1S $T=324260 678840 1 180 $X=323020 $Y=678460
X94 1770 2 1802 1 INV1S $T=325500 588120 1 180 $X=324260 $Y=587740
X95 1772 2 1796 1 INV1S $T=325500 608280 0 180 $X=324260 $Y=602860
X96 1762 2 1804 1 INV1S $T=327980 598200 1 180 $X=326740 $Y=597820
X97 1797 2 1818 1 INV1S $T=326740 688920 0 0 $X=326740 $Y=688540
X98 1816 2 1729 1 INV1S $T=327980 557880 1 0 $X=327980 $Y=552460
X99 124 2 1826 1 INV1S $T=329840 648600 1 180 $X=328600 $Y=648220
X100 1835 2 1661 1 INV1S $T=330460 678840 1 180 $X=329220 $Y=678460
X101 138 2 1847 1 INV1S $T=331080 658680 1 0 $X=331080 $Y=653260
X102 141 2 1815 1 INV1S $T=337280 638520 0 180 $X=336040 $Y=633100
X103 1864 2 1656 1 INV1S $T=336660 668760 0 0 $X=336660 $Y=668380
X104 1870 2 1876 1 INV1S $T=340380 567960 1 0 $X=340380 $Y=562540
X105 1863 2 1880 1 INV1S $T=341000 588120 0 0 $X=341000 $Y=587740
X106 1649 2 1593 1 INV1S $T=342860 588120 0 0 $X=342860 $Y=587740
X107 1869 2 1873 1 INV1S $T=344720 688920 0 180 $X=343480 $Y=683500
X108 1916 2 1885 1 INV1S $T=346580 688920 0 180 $X=345340 $Y=683500
X109 1864 2 1712 1 INV1S $T=347200 618360 0 180 $X=345960 $Y=612940
X110 1937 2 1886 1 INV1S $T=348440 567960 0 180 $X=347200 $Y=562540
X111 1945 2 1758 1 INV1S $T=350300 618360 0 180 $X=349060 $Y=612940
X112 1945 2 1629 1 INV1S $T=350300 668760 1 180 $X=349060 $Y=668380
X113 152 2 1934 1 INV1S $T=351540 648600 0 180 $X=350300 $Y=643180
X114 1871 2 1904 1 INV1S $T=350920 578040 0 0 $X=350920 $Y=577660
X115 165 2 1946 1 INV1S $T=352160 628440 1 180 $X=350920 $Y=628060
X116 159 2 1887 1 INV1S $T=352160 638520 0 180 $X=350920 $Y=633100
X117 1950 2 1931 1 INV1S $T=352780 588120 1 180 $X=351540 $Y=587740
X118 157 2 1881 1 INV1S $T=352780 638520 1 180 $X=351540 $Y=638140
X119 1775 2 1955 1 INV1S $T=352160 648600 1 0 $X=352160 $Y=643180
X120 1904 2 1950 1 INV1S $T=352780 578040 0 0 $X=352780 $Y=577660
X121 1955 2 1961 1 INV1S $T=353400 638520 0 0 $X=353400 $Y=638140
X122 171 2 1922 1 INV1S $T=355260 688920 1 180 $X=354020 $Y=688540
X123 1955 2 1966 1 INV1S $T=354640 648600 1 0 $X=354640 $Y=643180
X124 1971 2 1896 1 INV1S $T=356500 678840 0 180 $X=355260 $Y=673420
X125 160 2 174 1 INV1S $T=356500 678840 1 0 $X=356500 $Y=673420
X126 1969 2 1956 1 INV1S $T=358360 588120 1 180 $X=357120 $Y=587740
X127 1974 2 1893 1 INV1S $T=358980 547800 1 180 $X=357740 $Y=547420
X128 1922 2 177 1 INV1S $T=358980 668760 1 0 $X=358980 $Y=663340
X129 1979 2 1971 1 INV1S $T=359600 678840 1 0 $X=359600 $Y=673420
X130 1986 2 1908 1 INV1S $T=361460 567960 0 0 $X=361460 $Y=567580
X131 1997 2 1992 1 INV1S $T=363940 588120 1 180 $X=362700 $Y=587740
X132 2019 2 1935 1 INV1S $T=367660 668760 0 180 $X=366420 $Y=663340
X133 2018 2 2020 1 INV1S $T=366420 688920 1 0 $X=366420 $Y=683500
X134 153 2 187 1 INV1S $T=367660 668760 1 0 $X=367660 $Y=663340
X135 2032 2 1999 1 INV1S $T=368900 688920 0 180 $X=367660 $Y=683500
X136 2045 2 2008 1 INV1S $T=371380 678840 0 180 $X=370140 $Y=673420
X137 2049 2 1995 1 INV1S $T=372000 578040 0 180 $X=370760 $Y=572620
X138 2052 2 1919 1 INV1S $T=372620 557880 1 180 $X=371380 $Y=557500
X139 1995 2 2052 1 INV1S $T=372000 567960 0 0 $X=372000 $Y=567580
X140 2066 2 2053 1 INV1S $T=375100 598200 0 180 $X=373860 $Y=592780
X141 1904 2 2071 1 INV1S $T=376960 557880 0 0 $X=376960 $Y=557500
X142 1991 2 2089 1 INV1S $T=376960 688920 1 0 $X=376960 $Y=683500
X143 2058 2 2044 1 INV1S $T=377580 668760 0 0 $X=377580 $Y=668380
X144 1997 2 2100 1 INV1S $T=379440 578040 1 0 $X=379440 $Y=572620
X145 196 2 2106 1 INV1S $T=382540 588120 1 0 $X=382540 $Y=582700
X146 2107 2 2078 1 INV1S $T=383780 658680 1 180 $X=382540 $Y=658300
X147 2134 2 2056 1 INV1S $T=386260 628440 1 180 $X=385020 $Y=628060
X148 2131 2 2108 1 INV1S $T=386260 678840 0 180 $X=385020 $Y=673420
X149 2052 2 2127 1 INV1S $T=388740 557880 1 180 $X=387500 $Y=557500
X150 201 2 2153 1 INV1S $T=391840 578040 1 180 $X=390600 $Y=577660
X151 2148 2 2134 1 INV1S $T=390600 618360 1 0 $X=390600 $Y=612940
X152 2052 2 2162 1 INV1S $T=391840 557880 0 0 $X=391840 $Y=557500
X153 2134 2 2163 1 INV1S $T=391840 628440 0 0 $X=391840 $Y=628060
X154 2194 2 2164 1 INV1S $T=398040 658680 0 180 $X=396800 $Y=653260
X155 2195 2 2154 1 INV1S $T=399280 658680 1 180 $X=398040 $Y=658300
X156 2090 2 2207 1 INV1S $T=399900 578040 0 0 $X=399900 $Y=577660
X157 2135 2 2209 1 INV1S $T=399900 658680 0 0 $X=399900 $Y=658300
X158 2186 2 2221 1 INV1S $T=401760 658680 0 0 $X=401760 $Y=658300
X159 103 2 126 1 INV1S $T=404240 547800 1 0 $X=404240 $Y=542380
X160 165 2 214 1 INV1S $T=406100 537720 0 0 $X=406100 $Y=537340
X161 2179 2 2177 1 INV1S $T=406100 668760 1 0 $X=406100 $Y=663340
X162 210 2 2240 1 INV1S $T=407960 588120 0 180 $X=406720 $Y=582700
X163 2129 2 2268 1 INV1S $T=410440 648600 1 0 $X=410440 $Y=643180
X164 2173 2 2269 1 INV1S $T=411060 658680 1 0 $X=411060 $Y=653260
X165 2274 2 2260 1 INV1S $T=413540 557880 1 180 $X=412300 $Y=557500
X166 2274 2 226 1 INV1S $T=414160 547800 1 180 $X=412920 $Y=547420
X167 1925 2 216 1 INV1S $T=415400 557880 1 180 $X=414160 $Y=557500
X168 2014 2 232 1 INV1S $T=416640 578040 1 0 $X=416640 $Y=572620
X169 221 2 2274 1 INV1S $T=418500 547800 1 180 $X=417260 $Y=547420
X170 2252 2 2288 1 INV1S $T=417260 668760 0 0 $X=417260 $Y=668380
X171 2325 2 2181 1 INV1S $T=421600 688920 1 180 $X=420360 $Y=688540
X172 2305 2 2329 1 INV1S $T=421600 648600 0 0 $X=421600 $Y=648220
X173 2325 2 2265 1 INV1S $T=422840 699000 0 180 $X=421600 $Y=693580
X174 2345 2 2196 1 INV1S $T=425320 678840 0 180 $X=424080 $Y=673420
X175 2345 2 2294 1 INV1S $T=425320 678840 1 180 $X=424080 $Y=678460
X176 2334 2 2346 1 INV1S $T=425320 638520 0 0 $X=425320 $Y=638140
X177 2362 2 2369 1 INV1S $T=426560 567960 0 0 $X=426560 $Y=567580
X178 2243 2 2373 1 INV1S $T=427180 648600 0 0 $X=427180 $Y=648220
X179 2393 2 2405 1 INV1S $T=430900 557880 0 0 $X=430900 $Y=557500
X180 2400 2 2397 1 INV1S $T=433380 567960 0 180 $X=432140 $Y=562540
X181 2370 2 2396 1 INV1S $T=434000 638520 0 180 $X=432760 $Y=633100
X182 2404 2 2190 1 INV1S $T=434620 588120 1 180 $X=433380 $Y=587740
X183 2410 2 2404 1 INV1S $T=435860 588120 1 180 $X=434620 $Y=587740
X184 2404 2 2385 1 INV1S $T=434620 598200 1 0 $X=434620 $Y=592780
X185 1531 2 2418 1 INV1S $T=435860 618360 1 0 $X=435860 $Y=612940
X186 1842 2 2419 1 INV1S $T=435860 638520 0 0 $X=435860 $Y=638140
X187 2420 2 2325 1 INV1S $T=437100 658680 1 180 $X=435860 $Y=658300
X188 2133 2 2431 1 INV1S $T=436480 608280 1 0 $X=436480 $Y=602860
X189 2271 2 2428 1 INV1S $T=437720 618360 1 0 $X=437720 $Y=612940
X190 2388 2 2435 1 INV1S $T=437720 638520 0 0 $X=437720 $Y=638140
X191 2216 2 2444 1 INV1S $T=441440 588120 1 180 $X=440200 $Y=587740
X192 2453 2 2447 1 INV1S $T=444540 547800 1 180 $X=443300 $Y=547420
X193 2387 2 2401 1 INV1S $T=443300 648600 1 0 $X=443300 $Y=643180
X194 2350 2 2483 1 INV1S $T=447640 598200 1 180 $X=446400 $Y=597820
X195 2351 2 2466 1 INV1S $T=447640 608280 1 180 $X=446400 $Y=607900
X196 1576 2 2473 1 INV1S $T=447640 618360 1 180 $X=446400 $Y=617980
X197 260 2 2386 1 INV1S $T=448260 567960 1 180 $X=447020 $Y=567580
X198 1738 2 2506 1 INV1S $T=450120 628440 0 0 $X=450120 $Y=628060
X199 2501 2 2492 1 INV1S $T=450120 638520 1 0 $X=450120 $Y=633100
X200 2356 2 2508 1 INV1S $T=450740 648600 0 0 $X=450740 $Y=648220
X201 2504 2 2491 1 INV1S $T=455080 598200 1 180 $X=453840 $Y=597820
X202 2500 2 2512 1 INV1S $T=453840 608280 0 0 $X=453840 $Y=607900
X203 2172 2 2530 1 INV1S $T=455080 598200 0 0 $X=455080 $Y=597820
X204 2513 2 2507 1 INV1S $T=455700 588120 1 0 $X=455700 $Y=582700
X205 1840 2 2535 1 INV1S $T=455700 618360 0 0 $X=455700 $Y=617980
X206 1799 2 2587 1 INV1S $T=455700 628440 1 0 $X=455700 $Y=623020
X207 2389 2 2541 1 INV1S $T=458180 648600 0 180 $X=456940 $Y=643180
X208 2507 2 2555 1 INV1S $T=458180 588120 0 0 $X=458180 $Y=587740
X209 2016 2 2560 1 INV1S $T=458180 608280 0 0 $X=458180 $Y=607900
X210 2555 2 2504 1 INV1S $T=458800 598200 1 0 $X=458800 $Y=592780
X211 2431 2 2573 1 INV1S $T=460040 608280 1 0 $X=460040 $Y=602860
X212 2413 2 2540 1 INV1S $T=462520 638520 0 0 $X=462520 $Y=638140
X213 2236 2 2599 1 INV1S $T=465620 598200 1 0 $X=465620 $Y=592780
X214 2605 2 283 1 INV1S $T=467480 719160 1 180 $X=466240 $Y=718780
X215 2614 2 2460 1 INV1S $T=469340 598200 0 180 $X=468100 $Y=592780
X216 2081 2 2622 1 INV1S $T=469960 618360 1 0 $X=469960 $Y=612940
X217 2597 2 2680 1 INV1S $T=469960 628440 1 0 $X=469960 $Y=623020
X218 2633 2 2345 1 INV1S $T=473060 588120 1 180 $X=471820 $Y=587740
X219 2646 2 2577 1 INV1S $T=475540 578040 0 180 $X=474300 $Y=572620
X220 2659 2 276 1 INV1S $T=477400 557880 0 180 $X=476160 $Y=552460
X221 295 2 273 1 INV1S $T=477400 588120 1 180 $X=476160 $Y=587740
X222 2257 2 2660 1 INV1S $T=478640 608280 1 0 $X=478640 $Y=602860
X223 2672 2 2644 1 INV1S $T=480500 628440 0 0 $X=480500 $Y=628060
X224 2659 2 2678 1 INV1S $T=481120 567960 1 0 $X=481120 $Y=562540
X225 2709 2 2605 1 INV1S $T=486700 628440 1 180 $X=485460 $Y=628060
X226 312 2 2659 1 INV1S $T=487320 557880 1 180 $X=486080 $Y=557500
X227 315 2 2698 1 INV1S $T=488560 557880 1 180 $X=487320 $Y=557500
X228 316 2 2613 1 INV1S $T=488560 578040 0 180 $X=487320 $Y=572620
X229 2709 2 2713 1 INV1S $T=487320 628440 0 0 $X=487320 $Y=628060
X230 2709 2 2712 1 INV1S $T=489180 608280 1 180 $X=487940 $Y=607900
X231 2709 2 2707 1 INV1S $T=489180 618360 0 180 $X=487940 $Y=612940
X232 2709 2 2750 1 INV1S $T=487940 618360 0 0 $X=487940 $Y=617980
X233 2687 2 2528 1 INV1S $T=489180 588120 0 0 $X=489180 $Y=587740
X234 2630 2 2722 1 INV1S $T=491040 588120 0 180 $X=489800 $Y=582700
X235 322 2 2725 1 INV1S $T=492280 537720 1 180 $X=491040 $Y=537340
X236 2722 2 2728 1 INV1S $T=491660 588120 0 0 $X=491660 $Y=587740
X237 2709 2 2738 1 INV1S $T=491660 598200 1 0 $X=491660 $Y=592780
X238 323 2 254 1 INV1S $T=492900 608280 0 180 $X=491660 $Y=602860
X239 2630 2 2709 1 INV1S $T=494140 588120 0 0 $X=494140 $Y=587740
X240 2761 2 2758 1 INV1S $T=495380 658680 0 180 $X=494140 $Y=653260
X241 326 2 2782 1 INV1S $T=497240 547800 1 0 $X=497240 $Y=542380
X242 2761 2 2787 1 INV1S $T=501580 658680 1 180 $X=500340 $Y=658300
X243 2766 2 2761 1 INV1S $T=502820 658680 0 180 $X=501580 $Y=653260
X244 2573 2 2824 1 INV1S $T=504060 608280 1 0 $X=504060 $Y=602860
X245 338 2 2802 1 INV1S $T=505920 547800 0 180 $X=504680 $Y=542380
X246 363 2 2876 1 INV1S $T=517080 537720 1 180 $X=515840 $Y=537340
X247 364 2 2789 1 INV1S $T=517080 547800 1 180 $X=515840 $Y=547420
X248 369 2 2834 1 INV1S $T=520180 547800 0 180 $X=518940 $Y=542380
X249 2937 2 373 1 INV1S $T=525760 547800 0 180 $X=524520 $Y=542380
X250 378 2 2894 1 INV1S $T=526380 567960 1 180 $X=525140 $Y=567580
X251 2942 2 379 1 INV1S $T=528240 537720 1 180 $X=527000 $Y=537340
X252 377 2 2619 1 INV1S $T=527000 547800 1 0 $X=527000 $Y=542380
X253 380 2 2611 1 INV1S $T=528860 557880 0 180 $X=527620 $Y=552460
X254 2977 2 2981 1 INV1S $T=533200 658680 1 0 $X=533200 $Y=653260
X255 2932 2 2977 1 INV1S $T=533820 648600 1 0 $X=533820 $Y=643180
X256 3019 2 391 1 INV1S $T=536920 547800 0 180 $X=535680 $Y=542380
X257 2977 2 3010 1 INV1S $T=537540 648600 0 0 $X=537540 $Y=648220
X258 3024 2 2646 1 INV1S $T=540640 578040 0 0 $X=540640 $Y=577660
X259 3025 2 3006 1 INV1S $T=541880 638520 1 180 $X=540640 $Y=638140
X260 2764 2 3028 1 INV1S $T=544360 588120 1 0 $X=544360 $Y=582700
X261 3038 2 2612 1 INV1S $T=546220 567960 0 180 $X=544980 $Y=562540
X262 408 2 3048 1 INV1S $T=545600 719160 0 0 $X=545600 $Y=718780
X263 346 2 3070 1 INV1S $T=547460 578040 0 0 $X=547460 $Y=577660
X264 3060 2 2875 1 INV1S $T=548700 709080 1 180 $X=547460 $Y=708700
X265 415 2 2727 1 INV1S $T=549320 567960 0 180 $X=548080 $Y=562540
X266 393 2 418 1 INV1S $T=551800 537720 0 0 $X=551800 $Y=537340
X267 2824 2 3032 1 INV1S $T=554900 608280 1 0 $X=554900 $Y=602860
X268 331 2 426 1 INV1S $T=555520 547800 1 0 $X=555520 $Y=542380
X269 3120 2 2839 1 INV1S $T=561100 719160 0 180 $X=559860 $Y=713740
X270 432 2 3120 1 INV1S $T=561100 719160 1 0 $X=561100 $Y=713740
X271 3120 2 3132 1 INV1S $T=561720 709080 0 0 $X=561720 $Y=708700
X272 3060 2 3082 1 INV1S $T=562960 719160 1 0 $X=562960 $Y=713740
X273 3148 2 3004 1 INV1S $T=567300 628440 0 180 $X=566060 $Y=623020
X274 3166 2 3156 1 INV1S $T=569780 638520 0 0 $X=569780 $Y=638140
X275 2824 2 3219 1 INV1S $T=580320 608280 1 0 $X=580320 $Y=602860
X276 2824 2 3188 1 INV1S $T=580320 608280 0 0 $X=580320 $Y=607900
X277 484 2 3060 1 INV1S $T=581560 719160 0 180 $X=580320 $Y=713740
X278 3060 2 3246 1 INV1S $T=583420 709080 0 0 $X=583420 $Y=708700
X279 3237 2 3239 1 INV1S $T=589620 648600 1 180 $X=588380 $Y=648220
X280 3192 2 3207 1 INV1S $T=593960 608280 0 180 $X=592720 $Y=602860
X281 3342 2 3394 1 INV1S $T=613800 628440 0 0 $X=613800 $Y=628060
X282 3394 2 3356 1 INV1S $T=616900 618360 0 180 $X=615660 $Y=612940
X283 3413 2 3395 1 INV1S $T=618140 678840 1 0 $X=618140 $Y=673420
X284 3394 2 589 1 INV1S $T=623720 608280 0 0 $X=623720 $Y=607900
X285 596 2 3458 1 INV1S $T=625580 688920 1 0 $X=625580 $Y=683500
X286 3466 2 3342 1 INV1S $T=627440 678840 1 180 $X=626200 $Y=678460
X287 3452 2 593 1 INV1S $T=626200 688920 0 0 $X=626200 $Y=688540
X288 3434 2 3469 1 INV1S $T=627440 699000 1 0 $X=627440 $Y=693580
X289 607 2 611 1 INV1S $T=631780 719160 0 0 $X=631780 $Y=718780
X290 3048 2 620 1 INV1S $T=634260 719160 0 0 $X=634260 $Y=718780
X291 3510 2 3505 1 INV1S $T=635500 688920 0 0 $X=635500 $Y=688540
X292 3432 2 3530 1 INV1S $T=635500 709080 1 0 $X=635500 $Y=703660
X293 608 2 3537 1 INV1S $T=636740 628440 0 0 $X=636740 $Y=628060
X294 3540 2 3373 1 INV1S $T=638600 638520 1 180 $X=637360 $Y=638140
X295 499 2 3544 1 INV1S $T=638600 709080 1 0 $X=638600 $Y=703660
X296 3540 2 3518 1 INV1S $T=641080 638520 1 180 $X=639840 $Y=638140
X297 3571 2 628 1 INV1S $T=642940 719160 0 180 $X=641700 $Y=713740
X298 631 2 3541 1 INV1S $T=644180 699000 1 180 $X=642940 $Y=698620
X299 3540 2 3575 1 INV1S $T=643560 638520 1 0 $X=643560 $Y=633100
X300 3579 2 3573 1 INV1S $T=646660 699000 1 180 $X=645420 $Y=698620
X301 3626 2 3540 1 INV1S $T=656580 638520 0 0 $X=656580 $Y=638140
X302 648 2 652 1 INV1S $T=657200 547800 0 0 $X=657200 $Y=547420
X303 3658 2 3627 1 INV1S $T=659680 638520 1 180 $X=658440 $Y=638140
X304 3540 2 3659 1 INV1S $T=658440 648600 1 0 $X=658440 $Y=643180
X305 3615 2 3687 1 INV1S $T=663400 608280 1 0 $X=663400 $Y=602860
X306 3692 2 629 1 INV1S $T=665260 588120 1 180 $X=664020 $Y=587740
X307 658 2 3692 1 INV1S $T=665260 709080 1 0 $X=665260 $Y=703660
X308 3680 2 3707 1 INV1S $T=667120 557880 1 0 $X=667120 $Y=552460
X309 613 2 3726 1 INV1S $T=672080 699000 1 180 $X=670840 $Y=698620
X310 3701 2 3724 1 INV1S $T=673940 638520 1 0 $X=673940 $Y=633100
X311 3750 2 3791 1 INV1S $T=683240 608280 1 0 $X=683240 $Y=602860
X312 3791 2 3757 1 INV1S $T=683860 598200 1 0 $X=683860 $Y=592780
X313 3603 2 3798 1 INV1S $T=684480 588120 0 0 $X=684480 $Y=587740
X314 3791 2 3769 1 INV1S $T=684480 598200 0 0 $X=684480 $Y=597820
X315 3692 2 3822 1 INV1S $T=689440 618360 1 0 $X=689440 $Y=612940
X316 3798 2 693 1 INV1S $T=690680 578040 0 0 $X=690680 $Y=577660
X317 3798 2 3826 1 INV1S $T=691300 588120 1 0 $X=691300 $Y=582700
X318 3822 2 3845 1 INV1S $T=691300 618360 1 0 $X=691300 $Y=612940
X319 3692 2 3626 1 INV1S $T=693160 648600 0 180 $X=691920 $Y=643180
X320 3845 2 3750 1 INV1S $T=693780 618360 1 0 $X=693780 $Y=612940
X321 3832 2 3870 1 INV1S $T=695640 628440 1 0 $X=695640 $Y=623020
X322 3870 2 3624 1 INV1S $T=699980 598200 1 180 $X=698740 $Y=597820
X323 3859 2 3892 1 INV1S $T=700600 567960 0 0 $X=700600 $Y=567580
X324 3870 2 3888 1 INV1S $T=700600 598200 0 0 $X=700600 $Y=597820
X325 3692 2 3880 1 INV1S $T=704320 709080 1 0 $X=704320 $Y=703660
X326 3845 2 3914 1 INV1S $T=706180 608280 0 0 $X=706180 $Y=607900
X327 3892 2 3903 1 INV1S $T=709280 567960 0 0 $X=709280 $Y=567580
X328 3941 2 3876 1 INV1S $T=714240 557880 1 180 $X=713000 $Y=557500
X329 3769 2 3941 1 INV1S $T=714240 567960 0 0 $X=714240 $Y=567580
X330 3941 2 3955 1 INV1S $T=716100 567960 0 0 $X=716100 $Y=567580
X331 722 2 3974 1 INV1S $T=720440 719160 1 0 $X=720440 $Y=713740
X332 3985 2 3856 1 INV1S $T=724160 598200 0 180 $X=722920 $Y=592780
X333 3984 2 718 1 INV1S $T=724780 719160 0 180 $X=723540 $Y=713740
X334 4007 2 3916 1 INV1S $T=727880 567960 1 180 $X=726640 $Y=567580
X335 3995 2 4005 1 INV1S $T=726640 719160 1 0 $X=726640 $Y=713740
X336 3847 2 4007 1 INV1S $T=729740 567960 1 180 $X=728500 $Y=567580
X337 4022 2 3847 1 INV1S $T=730360 578040 1 180 $X=729120 $Y=577660
X338 4013 2 3771 1 INV1S $T=730360 688920 1 180 $X=729120 $Y=688540
X339 4021 2 3862 1 INV1S $T=731600 628440 0 180 $X=730360 $Y=623020
X340 4034 2 3843 1 INV1S $T=732840 658680 0 180 $X=731600 $Y=653260
X341 4029 2 3890 1 INV1S $T=733460 628440 1 180 $X=732220 $Y=628060
X342 4030 2 3811 1 INV1S $T=733460 648600 0 180 $X=732220 $Y=643180
X343 4039 2 3968 1 INV1S $T=735320 608280 1 180 $X=734080 $Y=607900
X344 3902 2 3966 1 INV1S $T=735320 688920 0 0 $X=735320 $Y=688540
X345 4052 2 737 1 INV1S $T=737180 547800 1 180 $X=735940 $Y=547420
X346 4050 2 3776 1 INV1S $T=737180 588120 0 180 $X=735940 $Y=582700
X347 4053 2 3946 1 INV1S $T=737180 608280 0 180 $X=735940 $Y=602860
X348 4051 2 3885 1 INV1S $T=737180 618360 0 180 $X=735940 $Y=612940
X349 4055 2 3897 1 INV1S $T=737800 699000 1 180 $X=736560 $Y=698620
X350 4056 2 3918 1 INV1S $T=737800 719160 0 180 $X=736560 $Y=713740
X351 3562 2 4061 1 INV1S $T=737800 688920 1 0 $X=737800 $Y=683500
X352 4062 2 3760 1 INV1S $T=739040 688920 1 180 $X=737800 $Y=688540
X353 655 2 4067 1 INV1S $T=739660 678840 1 0 $X=739660 $Y=673420
X354 4072 2 3678 1 INV1S $T=740900 688920 1 180 $X=739660 $Y=688540
X355 4069 2 3792 1 INV1S $T=741520 588120 0 180 $X=740280 $Y=582700
X356 3966 2 4082 1 INV1S $T=741520 709080 0 0 $X=741520 $Y=708700
X357 4083 2 3644 1 INV1S $T=743380 678840 0 0 $X=743380 $Y=678460
X358 762 2 4046 1 INV1S $T=744000 618360 1 0 $X=744000 $Y=612940
X359 4091 2 4013 1 INV1S $T=744620 709080 0 0 $X=744620 $Y=708700
X360 4062 2 4106 1 INV1S $T=745860 608280 0 0 $X=745860 $Y=607900
X361 4110 2 739 1 INV1S $T=747720 719160 1 180 $X=746480 $Y=718780
X362 740 2 4145 1 INV1S $T=752680 699000 0 0 $X=752680 $Y=698620
X363 4145 2 4140 1 INV1S $T=755160 699000 0 0 $X=755160 $Y=698620
X364 4170 2 3660 1 INV1S $T=758260 678840 1 180 $X=757020 $Y=678460
X365 4156 2 4062 1 INV1S $T=757020 699000 0 0 $X=757020 $Y=698620
X366 3996 2 781 1 INV1S $T=758260 598200 1 0 $X=758260 $Y=592780
X367 4176 2 4170 1 INV1S $T=759500 678840 1 180 $X=758260 $Y=678460
X368 780 2 4129 1 INV1S $T=759500 719160 0 180 $X=758260 $Y=713740
X369 4194 2 4126 1 INV1S $T=762600 658680 0 180 $X=761360 $Y=653260
X370 4140 2 4194 1 INV1S $T=761360 668760 0 0 $X=761360 $Y=668380
X371 783 2 668 1 INV1S $T=763220 709080 1 180 $X=761980 $Y=708700
X372 4194 2 4133 1 INV1S $T=764460 658680 0 0 $X=764460 $Y=658300
X373 4233 2 785 1 INV1S $T=771280 578040 0 180 $X=770040 $Y=572620
X374 4062 2 4216 1 INV1S $T=770040 699000 0 0 $X=770040 $Y=698620
X375 4007 2 4240 1 INV1S $T=771280 578040 1 0 $X=771280 $Y=572620
X376 4067 2 796 1 INV1S $T=771900 678840 1 0 $X=771900 $Y=673420
X377 4233 2 4265 1 INV1S $T=780580 618360 1 0 $X=780580 $Y=612940
X378 4293 2 4115 1 INV1S $T=783060 578040 0 180 $X=781820 $Y=572620
X379 4233 2 4313 1 INV1S $T=785540 618360 1 0 $X=785540 $Y=612940
X380 4233 2 4325 1 INV1S $T=787400 628440 0 0 $X=787400 $Y=628060
X381 4233 2 4326 1 INV1S $T=787400 648600 1 0 $X=787400 $Y=643180
X382 814 2 812 1 INV1S $T=791740 578040 1 0 $X=791740 $Y=572620
X383 4360 2 4225 1 INV1S $T=796080 618360 1 180 $X=794840 $Y=617980
X384 4362 2 819 1 INV1S $T=796080 678840 0 0 $X=796080 $Y=678460
X385 4360 2 4278 1 INV1S $T=797940 618360 1 180 $X=796700 $Y=617980
X386 3284 2 4362 1 INV1S $T=796700 658680 1 0 $X=796700 $Y=653260
X387 4082 2 4333 1 INV1S $T=797320 719160 1 0 $X=797320 $Y=713740
X388 4385 2 4304 1 INV1S $T=800420 628440 1 180 $X=799180 $Y=628060
X389 4362 2 4357 1 INV1S $T=800420 648600 1 0 $X=800420 $Y=643180
X390 4398 2 823 1 INV1S $T=802280 678840 1 180 $X=801040 $Y=678460
X391 4402 2 824 1 INV1S $T=803520 678840 1 180 $X=802280 $Y=678460
X392 4222 2 4406 1 INV1S $T=803520 678840 0 0 $X=803520 $Y=678460
X393 4417 2 4360 1 INV1S $T=808480 618360 1 180 $X=807240 $Y=617980
X394 4385 2 4417 1 INV1S $T=807240 628440 1 0 $X=807240 $Y=623020
X395 4360 2 4431 1 INV1S $T=808480 618360 0 0 $X=808480 $Y=617980
X396 4082 2 4390 1 INV1S $T=814060 709080 1 180 $X=812820 $Y=708700
X397 4456 2 834 1 INV1S $T=815300 537720 0 0 $X=815300 $Y=537340
X398 4082 2 4481 1 INV1S $T=817780 709080 0 0 $X=817780 $Y=708700
X399 4492 2 4393 1 INV1S $T=821500 557880 1 180 $X=820260 $Y=557500
X400 4492 2 4420 1 INV1S $T=821500 567960 0 180 $X=820260 $Y=562540
X401 849 2 4476 1 INV1S $T=821500 709080 1 0 $X=821500 $Y=703660
X402 4499 2 4492 1 INV1S $T=823360 567960 0 180 $X=822120 $Y=562540
X403 4522 2 4479 1 INV1S $T=825840 709080 0 0 $X=825840 $Y=708700
X404 4540 2 4556 1 INV1S $T=828320 699000 1 0 $X=828320 $Y=693580
X405 4564 2 4487 1 INV1S $T=833280 588120 0 180 $X=832040 $Y=582700
X406 4487 2 4579 1 INV1S $T=834520 608280 0 0 $X=834520 $Y=607900
X407 4534 2 4590 1 INV1S $T=835760 598200 1 0 $X=835760 $Y=592780
X408 4585 2 4578 1 INV1S $T=837000 608280 0 180 $X=835760 $Y=602860
X409 871 2 4568 1 INV1S $T=837000 699000 1 180 $X=835760 $Y=698620
X410 4492 2 4601 1 INV1S $T=836380 557880 0 0 $X=836380 $Y=557500
X411 4594 2 4604 1 INV1S $T=841340 608280 1 0 $X=841340 $Y=602860
X412 4615 2 4494 1 INV1S $T=841960 688920 1 0 $X=841960 $Y=683500
X413 4595 2 4385 1 INV1S $T=845680 628440 1 0 $X=845680 $Y=623020
X414 4637 2 4650 1 INV1S $T=845680 668760 1 0 $X=845680 $Y=663340
X415 3902 2 4595 1 INV1S $T=848160 628440 0 180 $X=846920 $Y=623020
X416 4566 2 4663 1 INV1S $T=848160 668760 1 0 $X=848160 $Y=663340
X417 4663 2 892 1 INV1S $T=851880 608280 0 0 $X=851880 $Y=607900
X418 4385 2 4683 1 INV1S $T=851880 618360 0 0 $X=851880 $Y=617980
X419 4385 2 4689 1 INV1S $T=851880 628440 1 0 $X=851880 $Y=623020
X420 4663 2 4690 1 INV1S $T=852500 668760 0 0 $X=852500 $Y=668380
X421 4704 2 4654 1 INV1S $T=856220 648600 0 180 $X=854980 $Y=643180
X422 894 2 4719 1 INV1S $T=855600 709080 0 0 $X=855600 $Y=708700
X423 4714 2 4704 1 INV1S $T=857460 648600 0 180 $X=856220 $Y=643180
X424 4061 2 900 1 INV1S $T=856840 688920 1 0 $X=856840 $Y=683500
X425 4742 2 891 1 INV1S $T=861800 588120 0 0 $X=861800 $Y=587740
X426 4582 2 4745 1 INV1S $T=863040 628440 0 0 $X=863040 $Y=628060
X427 4761 2 901 1 INV1S $T=865520 578040 1 180 $X=864280 $Y=577660
X428 4718 2 4761 1 INV1S $T=864280 588120 0 0 $X=864280 $Y=587740
X429 4751 2 897 1 INV1S $T=864900 598200 1 0 $X=864900 $Y=592780
X430 4061 2 4767 1 INV1S $T=865520 658680 1 0 $X=865520 $Y=653260
X431 4809 2 4727 1 INV1S $T=877300 648600 1 180 $X=876060 $Y=648220
X432 4850 2 4805 1 INV1S $T=881640 699000 0 180 $X=880400 $Y=693580
X433 4848 2 4813 1 INV1S $T=881020 578040 0 0 $X=881020 $Y=577660
X434 4852 2 4799 1 INV1S $T=881640 628440 0 0 $X=881640 $Y=628060
X435 3902 2 4870 1 INV1S $T=883500 688920 0 0 $X=883500 $Y=688540
X436 4840 2 4599 1 INV1S $T=884740 618360 0 0 $X=884740 $Y=617980
X437 4579 2 4856 1 INV1S $T=886600 608280 1 180 $X=885360 $Y=607900
X438 4850 2 4883 1 INV1S $T=885360 688920 0 0 $X=885360 $Y=688540
X439 4870 2 4850 1 INV1S $T=885360 699000 1 0 $X=885360 $Y=693580
X440 4875 2 821 1 INV1S $T=885980 588120 1 0 $X=885980 $Y=582700
X441 4813 2 4887 1 INV1S $T=886600 567960 0 0 $X=886600 $Y=567580
X442 4878 2 4499 1 INV1S $T=887840 578040 1 180 $X=886600 $Y=577660
X443 4878 2 4820 1 INV1S $T=886600 588120 0 0 $X=886600 $Y=587740
X444 4579 2 4888 1 INV1S $T=886600 608280 0 0 $X=886600 $Y=607900
X445 4875 2 922 1 INV1S $T=889080 578040 0 0 $X=889080 $Y=577660
X446 4898 2 4877 1 INV1S $T=889080 588120 0 0 $X=889080 $Y=587740
X447 4568 2 4760 1 INV1S $T=892800 628440 0 0 $X=892800 $Y=628060
X448 4875 2 4950 1 INV1S $T=897760 688920 1 0 $X=897760 $Y=683500
X449 4942 2 4935 1 INV1S $T=900240 557880 1 0 $X=900240 $Y=552460
X450 4942 2 4819 1 INV1S $T=900860 567960 1 0 $X=900860 $Y=562540
X451 960 2 961 1 INV1S $T=905200 719160 0 0 $X=905200 $Y=718780
X452 4690 2 5011 1 INV1S $T=907060 678840 1 0 $X=907060 $Y=673420
X453 5069 2 4944 1 INV1S $T=918840 578040 0 180 $X=917600 $Y=572620
X454 5078 2 4913 1 INV1S $T=920700 628440 1 180 $X=919460 $Y=628060
X455 5082 2 5078 1 INV1S $T=921940 628440 0 180 $X=920700 $Y=623020
X456 5078 2 4974 1 INV1S $T=921940 628440 0 0 $X=921940 $Y=628060
X457 5100 2 5069 1 INV1S $T=923800 578040 1 180 $X=922560 $Y=577660
X458 5011 2 5102 1 INV1S $T=923180 678840 0 0 $X=923180 $Y=678460
X459 4884 2 5144 1 INV1S $T=929380 648600 1 0 $X=929380 $Y=643180
X460 4599 2 986 1 INV1S $T=930620 547800 1 0 $X=930620 $Y=542380
X461 5139 2 5153 1 INV1S $T=931860 588120 1 0 $X=931860 $Y=582700
X462 5171 2 5196 1 INV1S $T=939300 598200 0 0 $X=939300 $Y=597820
X463 5205 2 5133 1 INV1S $T=941780 668760 1 180 $X=940540 $Y=668380
X464 5035 2 5205 1 INV1S $T=941160 678840 1 0 $X=941160 $Y=673420
X465 5221 2 989 1 INV1S $T=944260 557880 1 0 $X=944260 $Y=552460
X466 5221 2 5137 1 INV1S $T=945500 567960 0 180 $X=944260 $Y=562540
X467 5201 2 5221 1 INV1S $T=944260 567960 0 0 $X=944260 $Y=567580
X468 5240 2 5261 1 INV1S $T=947980 638520 0 0 $X=947980 $Y=638140
X469 5205 2 5255 1 INV1S $T=948600 678840 1 0 $X=948600 $Y=673420
X470 5091 2 5266 1 INV1S $T=955420 608280 0 0 $X=955420 $Y=607900
X471 5295 2 4967 1 INV1S $T=957900 567960 0 180 $X=956660 $Y=562540
X472 4887 2 5284 1 INV1S $T=956660 578040 1 0 $X=956660 $Y=572620
X473 4887 2 5278 1 INV1S $T=958520 557880 0 0 $X=958520 $Y=557500
X474 910 2 5295 1 INV1S $T=967820 547800 0 0 $X=967820 $Y=547420
X475 5295 2 5303 1 INV1S $T=970300 547800 1 180 $X=969060 $Y=547420
X476 4878 2 5243 1 INV1S $T=972160 618360 0 0 $X=972160 $Y=617980
X477 4685 2 5350 1 INV1S $T=972780 638520 0 0 $X=972780 $Y=638140
X478 5243 2 5362 1 INV1S $T=974020 618360 0 0 $X=974020 $Y=617980
X479 5362 2 5277 1 INV1S $T=974640 628440 1 0 $X=974640 $Y=623020
X480 5360 2 5368 1 INV1S $T=974640 699000 1 0 $X=974640 $Y=693580
X481 5362 2 5271 1 INV1S $T=976500 618360 1 180 $X=975260 $Y=617980
X482 5369 2 5345 1 INV1S $T=976500 588120 1 0 $X=976500 $Y=582700
X483 5295 2 1033 1 INV1S $T=977740 547800 1 0 $X=977740 $Y=542380
X484 5362 2 5364 1 INV1S $T=977740 618360 0 0 $X=977740 $Y=617980
X485 5362 2 5388 1 INV1S $T=980220 618360 0 0 $X=980220 $Y=617980
X486 5372 2 5412 1 INV1S $T=982700 618360 0 0 $X=982700 $Y=617980
X487 5406 2 5375 1 INV1S $T=982700 658680 0 0 $X=982700 $Y=658300
X488 5379 2 5417 1 INV1S $T=983940 678840 0 0 $X=983940 $Y=678460
X489 5424 2 1042 1 INV1S $T=986420 557880 0 180 $X=985180 $Y=552460
X490 1042 2 5428 1 INV1S $T=985800 547800 0 0 $X=985800 $Y=547420
X491 5393 2 5420 1 INV1S $T=986420 588120 1 0 $X=986420 $Y=582700
X492 983 2 5440 1 INV1S $T=987040 719160 1 0 $X=987040 $Y=713740
X493 5341 2 1049 1 INV1S $T=987660 547800 0 0 $X=987660 $Y=547420
X494 1049 2 1059 1 INV1S $T=990140 537720 0 0 $X=990140 $Y=537340
X495 5453 2 5466 1 INV1S $T=990140 648600 0 0 $X=990140 $Y=648220
X496 5457 2 5408 1 INV1S $T=990760 578040 0 0 $X=990760 $Y=577660
X497 5441 2 5469 1 INV1S $T=991380 678840 0 0 $X=991380 $Y=678460
X498 5464 2 1066 1 INV1S $T=991380 719160 0 0 $X=991380 $Y=718780
X499 5470 2 5467 1 INV1S $T=992620 578040 0 0 $X=992620 $Y=577660
X500 5464 2 5386 1 INV1S $T=994480 719160 1 180 $X=993240 $Y=718780
X501 5474 2 5464 1 INV1S $T=995720 719160 0 180 $X=994480 $Y=713740
X502 5466 2 5499 1 INV1S $T=996340 648600 0 0 $X=996340 $Y=648220
X503 5498 2 5522 1 INV1S $T=1001300 588120 0 0 $X=1001300 $Y=587740
X504 5345 2 5541 1 INV1S $T=1002540 598200 1 0 $X=1002540 $Y=592780
X505 5521 2 5547 1 INV1S $T=1005020 588120 1 0 $X=1005020 $Y=582700
X506 5295 2 5574 1 INV1S $T=1008740 547800 0 0 $X=1008740 $Y=547420
X507 5539 2 5614 1 INV1S $T=1014940 588120 0 0 $X=1014940 $Y=587740
X508 5614 2 1091 1 INV1S $T=1016180 567960 0 0 $X=1016180 $Y=567580
X509 5295 2 5637 1 INV1S $T=1018660 537720 0 0 $X=1018660 $Y=537340
X510 5614 2 5619 1 INV1S $T=1018660 578040 1 0 $X=1018660 $Y=572620
X511 4878 2 5575 1 INV1S $T=1020520 588120 0 0 $X=1020520 $Y=587740
X512 5455 2 5652 1 INV1S $T=1020520 658680 0 0 $X=1020520 $Y=658300
X513 5543 2 1099 1 INV1S $T=1023000 537720 1 180 $X=1021760 $Y=537340
X514 5659 2 5517 1 INV1S $T=1023620 578040 0 180 $X=1022380 $Y=572620
X515 5541 2 5654 1 INV1S $T=1023620 598200 1 180 $X=1022380 $Y=597820
X516 5673 2 1104 1 INV1S $T=1026100 719160 1 180 $X=1024860 $Y=718780
X517 1107 2 5673 1 INV1S $T=1027340 719160 1 180 $X=1026100 $Y=718780
X518 5652 2 5681 1 INV1S $T=1026720 658680 0 0 $X=1026720 $Y=658300
X519 5673 2 5611 1 INV1S $T=1027960 719160 1 0 $X=1027960 $Y=713740
X520 5717 2 5720 1 INV1S $T=1034780 578040 1 0 $X=1034780 $Y=572620
X521 4878 2 5721 1 INV1S $T=1034780 588120 0 0 $X=1034780 $Y=587740
X522 5541 2 5826 1 INV1S $T=1053380 598200 1 0 $X=1053380 $Y=592780
X523 5440 2 5747 1 INV1S $T=1055860 709080 0 0 $X=1055860 $Y=708700
X524 5721 2 5925 1 INV1S $T=1071360 578040 0 0 $X=1071360 $Y=577660
X525 5440 2 5936 1 INV1S $T=1073840 709080 0 0 $X=1073840 $Y=708700
X526 5998 2 5857 1 INV1S $T=1087480 688920 1 180 $X=1086240 $Y=688540
X527 5998 2 6001 1 INV1S $T=1087480 688920 0 0 $X=1087480 $Y=688540
X528 5989 2 5998 1 INV1S $T=1089340 699000 0 180 $X=1088100 $Y=693580
X529 5975 2 6032 1 INV1S $T=1093060 638520 1 0 $X=1093060 $Y=633100
X530 6032 2 5962 1 INV1S $T=1095540 638520 0 180 $X=1094300 $Y=633100
X531 1142 2 6066 1 INV1S $T=1099260 668760 1 0 $X=1099260 $Y=663340
X532 6032 2 6025 1 INV1S $T=1099880 638520 1 0 $X=1099880 $Y=633100
X533 6066 2 6005 1 INV1S $T=1100500 648600 0 0 $X=1100500 $Y=648220
X534 6066 2 6077 1 INV1S $T=1101740 668760 1 0 $X=1101740 $Y=663340
X535 5717 2 1178 1 INV1S $T=1103600 557880 0 0 $X=1103600 $Y=557500
X536 1177 2 6110 1 INV1S $T=1104220 537720 0 0 $X=1104220 $Y=537340
X537 6146 2 6159 1 INV1S $T=1113520 547800 1 0 $X=1113520 $Y=542380
X538 6075 2 1190 1 INV1S $T=1126540 537720 0 0 $X=1126540 $Y=537340
X539 6184 2 6182 1 INV1S $T=1128400 588120 0 180 $X=1127160 $Y=582700
X540 6002 2 6184 1 INV1S $T=1127160 598200 1 0 $X=1127160 $Y=592780
X541 6184 2 6181 1 INV1S $T=1128400 598200 1 180 $X=1127160 $Y=597820
X542 1235 1 2 1259 BUF1S $T=220720 608280 0 0 $X=220720 $Y=607900
X543 1264 1 2 1268 BUF1S $T=227540 588120 1 180 $X=225060 $Y=587740
X544 1282 1 2 10 BUF1S $T=230020 578040 0 0 $X=230020 $Y=577660
X545 1249 1 2 1282 BUF1S $T=234980 628440 0 180 $X=232500 $Y=623020
X546 1259 1 2 13 BUF1S $T=235600 557880 0 180 $X=233120 $Y=552460
X547 1312 1 2 1284 BUF1S $T=233120 699000 1 0 $X=233120 $Y=693580
X548 26 1 2 1369 BUF1S $T=243040 537720 0 0 $X=243040 $Y=537340
X549 37 1 2 1288 BUF1S $T=246140 699000 1 180 $X=243660 $Y=698620
X550 1393 1 2 39 BUF1S $T=249860 699000 1 180 $X=247380 $Y=698620
X551 1438 1 2 1264 BUF1S $T=253580 578040 1 180 $X=251100 $Y=577660
X552 1428 1 2 1410 BUF1S $T=253580 628440 1 180 $X=251100 $Y=628060
X553 42 1 2 1437 BUF1S $T=251100 699000 0 0 $X=251100 $Y=698620
X554 1438 1 2 21 BUF1S $T=254820 557880 0 180 $X=252340 $Y=552460
X555 1443 1 2 1414 BUF1S $T=255440 608280 1 180 $X=252960 $Y=607900
X556 43 1 2 1449 BUF1S $T=253580 719160 0 0 $X=253580 $Y=718780
X557 1465 1 2 1387 BUF1S $T=258540 547800 1 0 $X=258540 $Y=542380
X558 59 1 2 1469 BUF1S $T=262260 537720 1 180 $X=259780 $Y=537340
X559 1249 1 2 1483 BUF1S $T=259780 638520 1 0 $X=259780 $Y=633100
X560 1454 1 2 1397 BUF1S $T=262260 648600 1 180 $X=259780 $Y=648220
X561 79 1 2 1425 BUF1S $T=262260 678840 1 180 $X=259780 $Y=678460
X562 1437 1 2 1408 BUF1S $T=260400 608280 1 0 $X=260400 $Y=602860
X563 1443 1 2 1441 BUF1S $T=261640 628440 0 0 $X=261640 $Y=628060
X564 1501 1 2 1424 BUF1S $T=265360 648600 1 180 $X=262880 $Y=648220
X565 52 1 2 1398 BUF1S $T=267840 658680 0 180 $X=265360 $Y=653260
X566 1441 1 2 67 BUF1S $T=268460 709080 0 0 $X=268460 $Y=708700
X567 1530 1 2 1438 BUF1S $T=272800 578040 1 180 $X=270320 $Y=577660
X568 1511 1 2 61 BUF1S $T=274660 547800 0 180 $X=272180 $Y=542380
X569 1556 1 2 1399 BUF1S $T=276520 688920 1 180 $X=274040 $Y=688540
X570 1557 1 2 1506 BUF1S $T=275900 628440 1 0 $X=275900 $Y=623020
X571 1566 1 2 1558 BUF1S $T=279620 598200 1 180 $X=277140 $Y=597820
X572 1483 1 2 1562 BUF1S $T=277140 638520 0 0 $X=277140 $Y=638140
X573 1418 1 2 1566 BUF1S $T=277760 638520 1 0 $X=277760 $Y=633100
X574 46 1 2 1592 BUF1S $T=280240 567960 0 0 $X=280240 $Y=567580
X575 26 1 2 1587 BUF1S $T=280860 547800 1 0 $X=280860 $Y=542380
X576 1585 1 2 37 BUF1S $T=284580 719160 0 180 $X=282100 $Y=713740
X577 1623 1 2 1508 BUF1S $T=286440 618360 1 180 $X=283960 $Y=617980
X578 1469 1 2 1612 BUF1S $T=284580 557880 0 0 $X=284580 $Y=557500
X579 1543 1 2 83 BUF1S $T=285820 699000 1 0 $X=285820 $Y=693580
X580 1497 1 2 88 BUF1S $T=286440 588120 1 0 $X=286440 $Y=582700
X581 1578 1 2 1620 BUF1S $T=286440 618360 1 0 $X=286440 $Y=612940
X582 84 1 2 1585 BUF1S $T=288920 719160 0 180 $X=286440 $Y=713740
X583 44 1 2 1611 BUF1S $T=287680 567960 1 0 $X=287680 $Y=562540
X584 1629 1 2 1393 BUF1S $T=290780 699000 0 180 $X=288300 $Y=693580
X585 89 1 2 92 BUF1S $T=290160 537720 0 0 $X=290160 $Y=537340
X586 1387 1 2 1638 BUF1S $T=290160 557880 0 0 $X=290160 $Y=557500
X587 1562 1 2 1649 BUF1S $T=290780 588120 1 0 $X=290780 $Y=582700
X588 1629 1 2 95 BUF1S $T=290780 699000 1 0 $X=290780 $Y=693580
X589 1651 1 2 52 BUF1S $T=296980 678840 1 180 $X=294500 $Y=678460
X590 1556 1 2 1692 BUF1S $T=300080 678840 0 0 $X=300080 $Y=678460
X591 1675 1 2 1705 BUF1S $T=303180 567960 1 0 $X=303180 $Y=562540
X592 1566 1 2 1731 BUF1S $T=307520 588120 0 0 $X=307520 $Y=587740
X593 1752 1 2 1652 BUF1S $T=313100 709080 1 180 $X=310620 $Y=708700
X594 1761 1 2 1653 BUF1S $T=315580 557880 1 180 $X=313100 $Y=557500
X595 1743 1 2 1648 BUF1S $T=318680 557880 1 180 $X=316200 $Y=557500
X596 1794 1 2 1752 BUF1S $T=320540 678840 1 180 $X=318060 $Y=678460
X597 1743 1 2 1795 BUF1S $T=318680 557880 0 0 $X=318680 $Y=557500
X598 1794 1 2 1695 BUF1S $T=322400 668760 1 180 $X=319920 $Y=668380
X599 1418 1 2 1817 BUF1S $T=327360 638520 1 0 $X=327360 $Y=633100
X600 1483 1 2 1852 BUF1S $T=332320 648600 0 0 $X=332320 $Y=648220
X601 1816 1 2 1858 BUF1S $T=333560 578040 0 0 $X=333560 $Y=577660
X602 1886 1 2 1742 BUF1S $T=341000 557880 0 180 $X=338520 $Y=552460
X603 1885 1 2 1484 BUF1S $T=342240 678840 1 180 $X=339760 $Y=678460
X604 1649 1 2 1920 BUF1S $T=344720 588120 0 0 $X=344720 $Y=587740
X605 1917 1 2 1536 BUF1S $T=347200 608280 1 180 $X=344720 $Y=607900
X606 1886 1 2 1975 BUF1S $T=355260 567960 1 0 $X=355260 $Y=562540
X607 1731 1 2 1987 BUF1S $T=358980 588120 0 0 $X=358980 $Y=587740
X608 179 1 2 1794 BUF1S $T=362700 668760 0 180 $X=360220 $Y=663340
X609 1966 1 2 1984 BUF1S $T=366420 628440 0 0 $X=366420 $Y=628060
X610 1908 1 2 2041 BUF1S $T=368280 557880 0 0 $X=368280 $Y=557500
X611 1978 1 2 2070 BUF1S $T=373240 547800 1 0 $X=373240 $Y=542380
X612 2071 1 2 1911 BUF1S $T=375720 557880 1 180 $X=373240 $Y=557500
X613 2065 1 2 1974 BUF1S $T=375720 567960 0 180 $X=373240 $Y=562540
X614 2071 1 2 2097 BUF1S $T=378820 557880 0 0 $X=378820 $Y=557500
X615 2100 1 2 1973 BUF1S $T=385020 567960 0 180 $X=382540 $Y=562540
X616 2121 1 2 197 BUF1S $T=385020 688920 0 180 $X=382540 $Y=683500
X617 203 1 2 200 BUF1S $T=386260 719160 1 180 $X=383780 $Y=718780
X618 2139 1 2 2051 BUF1S $T=389360 668760 0 180 $X=386880 $Y=663340
X619 1961 1 2 2123 BUF1S $T=387500 628440 0 0 $X=387500 $Y=628060
X620 2116 1 2 2009 BUF1S $T=389980 678840 0 180 $X=387500 $Y=673420
X621 2096 1 2 204 BUF1S $T=389980 709080 1 180 $X=387500 $Y=708700
X622 2143 1 2 199 BUF1S $T=389980 719160 1 180 $X=387500 $Y=718780
X623 1961 1 2 2112 BUF1S $T=389360 638520 1 0 $X=389360 $Y=633100
X624 2154 1 2 208 BUF1S $T=391220 678840 0 0 $X=391220 $Y=678460
X625 2208 1 2 1917 BUF1S $T=400520 598200 0 180 $X=398040 $Y=592780
X626 2039 1 2 2234 BUF1S $T=405480 557880 0 0 $X=405480 $Y=557500
X627 2123 1 2 2212 BUF1S $T=407340 618360 1 0 $X=407340 $Y=612940
X628 2112 1 2 2253 BUF1S $T=407340 648600 1 0 $X=407340 $Y=643180
X629 2254 1 2 2169 BUF1S $T=409820 719160 0 180 $X=407340 $Y=713740
X630 224 1 2 188 BUF1S $T=412920 709080 1 180 $X=410440 $Y=708700
X631 198 1 2 228 BUF1S $T=410440 719160 1 0 $X=410440 $Y=713740
X632 2143 1 2 225 BUF1S $T=410440 719160 0 0 $X=410440 $Y=718780
X633 2227 1 2 227 BUF1S $T=411060 688920 1 0 $X=411060 $Y=683500
X634 218 1 2 2256 BUF1S $T=414160 547800 0 0 $X=414160 $Y=547420
X635 2317 1 2 233 BUF1S $T=419740 688920 1 0 $X=419740 $Y=683500
X636 2298 1 2 2138 BUF1S $T=424080 638520 1 180 $X=421600 $Y=638140
X637 2301 1 2 2139 BUF1S $T=424080 658680 1 180 $X=421600 $Y=658300
X638 2346 1 2 229 BUF1S $T=425940 648600 1 180 $X=423460 $Y=648220
X639 2391 1 2 236 BUF1S $T=430900 658680 0 180 $X=428420 $Y=653260
X640 2342 1 2 242 BUF1S $T=432140 719160 0 180 $X=429660 $Y=713740
X641 2380 1 2 2208 BUF1S $T=433380 588120 1 180 $X=430900 $Y=587740
X642 2401 1 2 2116 BUF1S $T=434620 658680 1 180 $X=432140 $Y=658300
X643 2383 1 2 231 BUF1S $T=432760 719160 1 0 $X=432760 $Y=713740
X644 2414 1 2 2277 BUF1S $T=436480 648600 0 180 $X=434000 $Y=643180
X645 2436 1 2 2254 BUF1S $T=440200 688920 0 180 $X=437720 $Y=683500
X646 2387 1 2 2301 BUF1S $T=442060 648600 1 180 $X=439580 $Y=648220
X647 2460 1 2 198 BUF1S $T=443300 688920 0 180 $X=440820 $Y=683500
X648 2366 1 2 249 BUF1S $T=442680 678840 1 0 $X=442680 $Y=673420
X649 2474 1 2 2322 BUF1S $T=445780 648600 1 180 $X=443300 $Y=648220
X650 237 1 2 2479 BUF1S $T=446400 537720 0 0 $X=446400 $Y=537340
X651 2514 1 2 224 BUF1S $T=453220 709080 1 180 $X=450740 $Y=708700
X652 2504 1 2 2500 BUF1S $T=456320 618360 0 180 $X=453840 $Y=612940
X653 2513 1 2 2539 BUF1S $T=455080 608280 1 0 $X=455080 $Y=602860
X654 2528 1 2 183 BUF1S $T=455080 709080 0 0 $X=455080 $Y=708700
X655 2507 1 2 2547 BUF1S $T=455700 608280 0 0 $X=455700 $Y=607900
X656 2504 1 2 2481 BUF1S $T=456940 638520 1 0 $X=456940 $Y=633100
X657 273 1 2 2565 BUF1S $T=463140 557880 1 180 $X=460660 $Y=557500
X658 2577 1 2 2143 BUF1S $T=463140 588120 1 180 $X=460660 $Y=587740
X659 2528 1 2 280 BUF1S $T=462520 567960 1 0 $X=462520 $Y=562540
X660 2619 1 2 2259 BUF1S $T=469960 588120 1 180 $X=467480 $Y=587740
X661 2584 1 2 2383 BUF1S $T=471200 578040 0 180 $X=468720 $Y=572620
X662 298 1 2 2588 BUF1S $T=479880 547800 0 180 $X=477400 $Y=542380
X663 300 1 2 282 BUF1S $T=480500 557880 0 180 $X=478020 $Y=552460
X664 297 1 2 2671 BUF1S $T=478640 557880 0 0 $X=478640 $Y=557500
X665 2668 1 2 2641 BUF1S $T=484220 618360 1 180 $X=481740 $Y=617980
X666 2641 1 2 2664 BUF1S $T=483600 648600 1 0 $X=483600 $Y=643180
X667 273 1 2 2514 BUF1S $T=485460 618360 0 0 $X=485460 $Y=617980
X668 2688 1 2 2642 BUF1S $T=486700 658680 1 0 $X=486700 $Y=653260
X669 2727 1 2 2436 BUF1S $T=491040 578040 0 180 $X=488560 $Y=572620
X670 2583 1 2 2688 BUF1S $T=491660 628440 1 180 $X=489180 $Y=628060
X671 2764 1 2 2584 BUF1S $T=496000 547800 0 180 $X=493520 $Y=542380
X672 2729 1 2 2766 BUF1S $T=496000 608280 0 0 $X=496000 $Y=607900
X673 2789 1 2 2617 BUF1S $T=500340 547800 1 180 $X=497860 $Y=547420
X674 2793 1 2 2762 BUF1S $T=501580 668760 0 180 $X=499100 $Y=663340
X675 2802 1 2 2593 BUF1S $T=504060 547800 0 180 $X=501580 $Y=542380
X676 2573 1 2 2807 BUF1S $T=501580 628440 0 0 $X=501580 $Y=628060
X677 2775 1 2 2793 BUF1S $T=504680 628440 0 0 $X=504680 $Y=628060
X678 2741 1 2 2734 BUF1S $T=509020 678840 0 180 $X=506540 $Y=673420
X679 2894 1 2 2420 BUF1S $T=519560 578040 0 180 $X=517080 $Y=572620
X680 2920 1 2 2266 BUF1S $T=523280 578040 1 180 $X=520800 $Y=577660
X681 384 1 2 2788 BUF1S $T=529480 709080 1 180 $X=527000 $Y=708700
X682 2805 1 2 2991 BUF1S $T=534440 618360 0 0 $X=534440 $Y=617980
X683 2991 1 2 2959 BUF1S $T=535060 658680 0 0 $X=535060 $Y=658300
X684 3006 1 2 2887 BUF1S $T=539400 618360 1 180 $X=536920 $Y=617980
X685 378 1 2 399 BUF1S $T=538780 547800 1 0 $X=538780 $Y=542380
X686 3024 1 2 3025 BUF1S $T=540640 588120 1 0 $X=540640 $Y=582700
X687 406 1 2 2764 BUF1S $T=544360 578040 0 0 $X=544360 $Y=577660
X688 3006 1 2 3031 BUF1S $T=549940 658680 0 180 $X=547460 $Y=653260
X689 2651 1 2 3081 BUF1S $T=549320 648600 0 0 $X=549320 $Y=648220
X690 384 1 2 3017 BUF1S $T=549320 699000 0 0 $X=549320 $Y=698620
X691 3069 1 2 3085 BUF1S $T=550560 648600 1 0 $X=550560 $Y=643180
X692 420 1 2 3038 BUF1S $T=553660 567960 0 180 $X=551180 $Y=562540
X693 2680 1 2 3092 BUF1S $T=551180 658680 0 0 $X=551180 $Y=658300
X694 3042 1 2 3069 BUF1S $T=553040 628440 0 0 $X=553040 $Y=628060
X695 3033 1 2 3104 BUF1S $T=554900 638520 0 0 $X=554900 $Y=638140
X696 447 1 2 3096 BUF1S $T=564200 537720 1 180 $X=561720 $Y=537340
X697 2624 1 2 3150 BUF1S $T=565440 638520 1 0 $X=565440 $Y=633100
X698 452 1 2 2962 BUF1S $T=567920 719160 0 180 $X=565440 $Y=713740
X699 3017 1 2 3171 BUF1S $T=568540 678840 0 0 $X=568540 $Y=678460
X700 3207 1 2 3110 BUF1S $T=580320 618360 1 180 $X=577840 $Y=617980
X701 3218 1 2 3151 BUF1S $T=582800 588120 0 0 $X=582800 $Y=587740
X702 3234 1 2 3094 BUF1S $T=585280 628440 0 180 $X=582800 $Y=623020
X703 3107 1 2 3186 BUF1S $T=586520 618360 0 0 $X=586520 $Y=617980
X704 3242 1 2 3172 BUF1S $T=590240 598200 0 0 $X=590240 $Y=597820
X705 3295 1 2 3241 BUF1S $T=593340 648600 0 0 $X=593340 $Y=648220
X706 3275 1 2 3285 BUF1S $T=598300 709080 0 0 $X=598300 $Y=708700
X707 3303 1 2 3329 BUF1S $T=599540 618360 0 0 $X=599540 $Y=617980
X708 471 1 2 3321 BUF1S $T=602640 547800 0 0 $X=602640 $Y=547420
X709 3342 1 2 3265 BUF1S $T=605120 658680 1 180 $X=602640 $Y=658300
X710 544 1 2 3159 BUF1S $T=605120 719160 0 180 $X=602640 $Y=713740
X711 3243 1 2 3307 BUF1S $T=604500 668760 1 0 $X=604500 $Y=663340
X712 3310 1 2 3354 BUF1S $T=604500 678840 1 0 $X=604500 $Y=673420
X713 3307 1 2 549 BUF1S $T=610080 638520 1 0 $X=610080 $Y=633100
X714 3374 1 2 3369 BUF1S $T=610700 608280 1 0 $X=610700 $Y=602860
X715 3373 1 2 1967 BUF1S $T=613800 658680 0 180 $X=611320 $Y=653260
X716 3343 1 2 3434 BUF1S $T=621860 678840 0 0 $X=621860 $Y=678460
X717 3440 1 2 3404 BUF1S $T=624960 638520 1 0 $X=624960 $Y=633100
X718 602 1 2 3368 BUF1S $T=629920 719160 0 180 $X=627440 $Y=713740
X719 3469 1 2 3494 BUF1S $T=629300 699000 1 0 $X=629300 $Y=693580
X720 3373 1 2 3499 BUF1S $T=631160 638520 0 0 $X=631160 $Y=638140
X721 608 1 2 617 BUF1S $T=631780 628440 0 0 $X=631780 $Y=628060
X722 3499 1 2 3353 BUF1S $T=633020 598200 0 0 $X=633020 $Y=597820
X723 3518 1 2 3310 BUF1S $T=635500 668760 0 180 $X=633020 $Y=663340
X724 3541 1 2 3275 BUF1S $T=638600 699000 1 180 $X=636120 $Y=698620
X725 639 1 2 580 BUF1S $T=646660 719160 1 180 $X=644180 $Y=718780
X726 3587 1 2 602 BUF1S $T=648520 719160 0 180 $X=646040 $Y=713740
X727 2798 1 2 643 BUF1S $T=651620 578040 1 0 $X=651620 $Y=572620
X728 3627 1 2 646 BUF1S $T=656580 618360 1 180 $X=654100 $Y=617980
X729 3644 1 2 3553 BUF1S $T=658440 678840 1 180 $X=655960 $Y=678460
X730 3678 1 2 3585 BUF1S $T=663400 688920 1 180 $X=660920 $Y=688540
X731 3645 1 2 3561 BUF1S $T=664640 688920 0 0 $X=664640 $Y=688540
X732 656 1 2 3701 BUF1S $T=664640 699000 0 0 $X=664640 $Y=698620
X733 3681 1 2 660 BUF1S $T=665880 537720 0 0 $X=665880 $Y=537340
X734 3698 1 2 3709 BUF1S $T=670840 598200 1 0 $X=670840 $Y=592780
X735 3757 1 2 3680 BUF1S $T=674560 578040 0 180 $X=672080 $Y=572620
X736 3537 1 2 3768 BUF1S $T=675180 648600 1 0 $X=675180 $Y=643180
X737 674 1 2 3571 BUF1S $T=678900 709080 1 180 $X=676420 $Y=708700
X738 3776 1 2 3721 BUF1S $T=681380 578040 0 180 $X=678900 $Y=572620
X739 3724 1 2 679 BUF1S $T=680140 638520 1 0 $X=680140 $Y=633100
X740 3811 1 2 3693 BUF1S $T=688200 638520 1 180 $X=685720 $Y=638140
X741 3803 1 2 3747 BUF1S $T=688200 678840 1 180 $X=685720 $Y=678460
X742 3792 1 2 3741 BUF1S $T=686960 567960 1 0 $X=686960 $Y=562540
X743 3824 1 2 3694 BUF1S $T=690060 678840 0 180 $X=687580 $Y=673420
X744 3803 1 2 3645 BUF1S $T=690680 699000 1 180 $X=688200 $Y=698620
X745 3822 1 2 3700 BUF1S $T=689440 628440 1 0 $X=689440 $Y=623020
X746 3843 1 2 3702 BUF1S $T=693780 648600 1 180 $X=691300 $Y=648220
X747 701 1 2 667 BUF1S $T=695640 537720 1 180 $X=693160 $Y=537340
X748 3862 1 2 3752 BUF1S $T=697500 618360 1 180 $X=695020 $Y=617980
X749 3859 1 2 3723 BUF1S $T=698740 638520 1 180 $X=696260 $Y=638140
X750 3873 1 2 3742 BUF1S $T=700600 648600 0 180 $X=698120 $Y=643180
X751 3885 1 2 3695 BUF1S $T=701220 618360 1 180 $X=698740 $Y=617980
X752 3890 1 2 3630 BUF1S $T=703080 648600 0 180 $X=700600 $Y=643180
X753 3880 1 2 674 BUF1S $T=703080 719160 0 180 $X=700600 $Y=713740
X754 3700 1 2 3806 BUF1S $T=701840 618360 0 0 $X=701840 $Y=617980
X755 3897 1 2 3713 BUF1S $T=704320 699000 1 180 $X=701840 $Y=698620
X756 708 1 2 3774 BUF1S $T=708040 598200 1 180 $X=705560 $Y=597820
X757 3880 1 2 3803 BUF1S $T=708040 699000 1 180 $X=705560 $Y=698620
X758 3918 1 2 3732 BUF1S $T=709900 709080 0 180 $X=707420 $Y=703660
X759 3880 1 2 711 BUF1S $T=707420 719160 1 0 $X=707420 $Y=713740
X760 3944 1 2 3900 BUF1S $T=715480 678840 0 180 $X=713000 $Y=673420
X761 3946 1 2 3595 BUF1S $T=716100 598200 1 180 $X=713620 $Y=597820
X762 3856 1 2 3858 BUF1S $T=717960 557880 1 180 $X=715480 $Y=557500
X763 719 1 2 3587 BUF1S $T=717960 719160 0 180 $X=715480 $Y=713740
X764 3968 1 2 3567 BUF1S $T=721060 598200 1 180 $X=718580 $Y=597820
X765 3978 1 2 3725 BUF1S $T=722300 668760 0 0 $X=722300 $Y=668380
X766 3856 1 2 4020 BUF1S $T=727260 588120 0 0 $X=727260 $Y=587740
X767 3912 1 2 3986 BUF1S $T=728500 638520 0 0 $X=728500 $Y=638140
X768 4019 1 2 3730 BUF1S $T=731600 648600 1 180 $X=729120 $Y=648220
X769 3900 1 2 3912 BUF1S $T=731600 658680 0 180 $X=729120 $Y=653260
X770 3955 1 2 4026 BUF1S $T=730360 567960 0 0 $X=730360 $Y=567580
X771 3862 1 2 4041 BUF1S $T=731600 628440 1 0 $X=731600 $Y=623020
X772 4024 1 2 736 BUF1S $T=732220 547800 0 0 $X=732220 $Y=547420
X773 4026 1 2 4040 BUF1S $T=732220 557880 1 0 $X=732220 $Y=552460
X774 3776 1 2 4042 BUF1S $T=733460 578040 0 0 $X=733460 $Y=577660
X775 3968 1 2 4043 BUF1S $T=733460 608280 1 0 $X=733460 $Y=602860
X776 3843 1 2 4048 BUF1S $T=734080 658680 1 0 $X=734080 $Y=653260
X777 740 1 2 3944 BUF1S $T=736560 699000 1 180 $X=734080 $Y=698620
X778 739 1 2 743 BUF1S $T=735320 628440 0 0 $X=735320 $Y=628060
X779 745 1 2 4060 BUF1S $T=737800 608280 0 0 $X=737800 $Y=607900
X780 749 1 2 753 BUF1S $T=737800 628440 0 0 $X=737800 $Y=628060
X781 3918 1 2 4066 BUF1S $T=737800 699000 0 0 $X=737800 $Y=698620
X782 3678 1 2 4076 BUF1S $T=739660 688920 1 0 $X=739660 $Y=683500
X783 4049 1 2 4024 BUF1S $T=742140 699000 0 180 $X=739660 $Y=693580
X784 3885 1 2 4079 BUF1S $T=740900 618360 1 0 $X=740900 $Y=612940
X785 764 1 2 756 BUF1S $T=743380 628440 1 180 $X=740900 $Y=628060
X786 760 1 2 744 BUF1S $T=743380 638520 0 180 $X=740900 $Y=633100
X787 757 1 2 4077 BUF1S $T=740900 699000 0 0 $X=740900 $Y=698620
X788 3897 1 2 4090 BUF1S $T=742140 699000 1 0 $X=742140 $Y=693580
X789 3946 1 2 4095 BUF1S $T=742760 608280 0 0 $X=742760 $Y=607900
X790 3890 1 2 4104 BUF1S $T=744000 638520 1 0 $X=744000 $Y=633100
X791 3644 1 2 4108 BUF1S $T=744620 688920 1 0 $X=744620 $Y=683500
X792 766 1 2 4027 BUF1S $T=747100 699000 0 180 $X=744620 $Y=693580
X793 732 1 2 4134 BUF1S $T=750200 547800 0 0 $X=750200 $Y=547420
X794 3811 1 2 4153 BUF1S $T=753920 648600 1 0 $X=753920 $Y=643180
X795 663 1 2 4107 BUF1S $T=755160 699000 1 0 $X=755160 $Y=693580
X796 3610 1 2 783 BUF1S $T=758880 709080 0 0 $X=758880 $Y=708700
X797 748 1 2 4183 BUF1S $T=764460 598200 0 180 $X=761980 $Y=592780
X798 4133 1 2 4217 BUF1S $T=765700 658680 0 0 $X=765700 $Y=658300
X799 787 1 2 4252 BUF1S $T=771900 699000 0 0 $X=771900 $Y=698620
X800 4180 1 2 4260 BUF1S $T=775000 678840 0 0 $X=775000 $Y=678460
X801 4148 1 2 4283 BUF1S $T=778100 648600 1 0 $X=778100 $Y=643180
X802 4365 1 2 4220 BUF1S $T=798560 557880 0 180 $X=796080 $Y=552460
X803 4352 1 2 4378 BUF1S $T=796080 709080 0 0 $X=796080 $Y=708700
X804 807 1 2 4210 BUF1S $T=796700 688920 1 0 $X=796700 $Y=683500
X805 4365 1 2 811 BUF1S $T=802280 557880 0 180 $X=799800 $Y=552460
X806 821 1 2 4396 BUF1S $T=800420 567960 1 0 $X=800420 $Y=562540
X807 4396 1 2 4144 BUF1S $T=804140 557880 1 180 $X=801660 $Y=557500
X808 4420 1 2 4365 BUF1S $T=807240 557880 1 180 $X=804760 $Y=557500
X809 4462 1 2 4442 BUF1S $T=815300 709080 0 0 $X=815300 $Y=708700
X810 814 1 2 4456 BUF1S $T=816540 537720 0 0 $X=816540 $Y=537340
X811 4481 1 2 4446 BUF1S $T=820260 688920 1 180 $X=817780 $Y=688540
X812 851 1 2 4521 BUF1S $T=823980 709080 1 0 $X=823980 $Y=703660
X813 858 1 2 862 BUF1S $T=826460 628440 1 0 $X=826460 $Y=623020
X814 4479 1 2 4544 BUF1S $T=827080 709080 0 0 $X=827080 $Y=708700
X815 4393 1 2 847 BUF1S $T=830180 537720 1 180 $X=827700 $Y=537340
X816 4517 1 2 4495 BUF1S $T=828320 709080 1 0 $X=828320 $Y=703660
X817 4556 1 2 4486 BUF1S $T=830180 699000 1 0 $X=830180 $Y=693580
X818 821 1 2 4525 BUF1S $T=831420 578040 0 0 $X=831420 $Y=577660
X819 4562 1 2 4508 BUF1S $T=831420 648600 0 0 $X=831420 $Y=648220
X820 4578 1 2 4530 BUF1S $T=835760 598200 1 180 $X=833280 $Y=597820
X821 873 1 2 870 BUF1S $T=839480 557880 0 180 $X=837000 $Y=552460
X822 4577 1 2 866 BUF1S $T=837620 567960 0 0 $X=837620 $Y=567580
X823 4027 1 2 4617 BUF1S $T=838860 658680 1 0 $X=838860 $Y=653260
X824 822 1 2 4625 BUF1S $T=840720 557880 1 0 $X=840720 $Y=552460
X825 4609 1 2 879 BUF1S $T=840720 598200 1 0 $X=840720 $Y=592780
X826 4610 1 2 4550 BUF1S $T=844440 648600 1 180 $X=841960 $Y=648220
X827 863 1 2 868 BUF1S $T=845060 567960 1 180 $X=842580 $Y=567580
X828 884 1 2 881 BUF1S $T=845060 618360 1 180 $X=842580 $Y=617980
X829 4595 1 2 4458 BUF1S $T=845060 628440 0 180 $X=842580 $Y=623020
X830 4581 1 2 4627 BUF1S $T=843200 709080 1 0 $X=843200 $Y=703660
X831 4046 1 2 4652 BUF1S $T=843820 598200 1 0 $X=843820 $Y=592780
X832 4464 1 2 887 BUF1S $T=844440 719160 1 0 $X=844440 $Y=713740
X833 4562 1 2 4660 BUF1S $T=845680 658680 0 0 $X=845680 $Y=658300
X834 869 1 2 4658 BUF1S $T=846300 588120 0 0 $X=846300 $Y=587740
X835 878 1 2 890 BUF1S $T=849400 628440 1 0 $X=849400 $Y=623020
X836 4672 1 2 4610 BUF1S $T=851880 658680 0 180 $X=849400 $Y=653260
X837 4673 1 2 4528 BUF1S $T=851880 668760 1 180 $X=849400 $Y=668380
X838 4494 1 2 4701 BUF1S $T=851260 688920 1 0 $X=851260 $Y=683500
X839 887 1 2 4651 BUF1S $T=851260 709080 1 0 $X=851260 $Y=703660
X840 4689 1 2 4705 BUF1S $T=853120 628440 1 0 $X=853120 $Y=623020
X841 4697 1 2 4713 BUF1S $T=854980 638520 0 0 $X=854980 $Y=638140
X842 4544 1 2 4733 BUF1S $T=858080 709080 1 0 $X=858080 $Y=703660
X843 4486 1 2 4725 BUF1S $T=859940 699000 1 0 $X=859940 $Y=693580
X844 4760 1 2 4557 BUF1S $T=864280 658680 0 180 $X=861800 $Y=653260
X845 4673 1 2 4744 BUF1S $T=864280 678840 1 0 $X=864280 $Y=673420
X846 4500 1 2 4743 BUF1S $T=866760 638520 0 0 $X=866760 $Y=638140
X847 4709 1 2 4783 BUF1S $T=867380 688920 1 0 $X=867380 $Y=683500
X848 4820 1 2 907 BUF1S $T=877300 567960 1 180 $X=874820 $Y=567580
X849 4821 1 2 4827 BUF1S $T=876060 598200 1 0 $X=876060 $Y=592780
X850 4578 1 2 4831 BUF1S $T=876060 598200 0 0 $X=876060 $Y=597820
X851 4799 1 2 4731 BUF1S $T=879780 628440 1 180 $X=877300 $Y=628060
X852 4727 1 2 4822 BUF1S $T=877300 648600 0 0 $X=877300 $Y=648220
X853 4805 1 2 4738 BUF1S $T=880400 699000 0 180 $X=877920 $Y=693580
X854 4829 1 2 4855 BUF1S $T=879160 598200 0 0 $X=879160 $Y=597820
X855 810 1 2 928 BUF1S $T=879780 618360 0 0 $X=879780 $Y=617980
X856 4805 1 2 4778 BUF1S $T=880400 709080 0 0 $X=880400 $Y=708700
X857 4736 1 2 4668 BUF1S $T=882260 618360 0 0 $X=882260 $Y=617980
X858 4877 1 2 913 BUF1S $T=885980 588120 1 180 $X=883500 $Y=587740
X859 4859 1 2 4871 BUF1S $T=884120 658680 1 0 $X=884120 $Y=653260
X860 4846 1 2 4896 BUF1S $T=885980 688920 1 0 $X=885980 $Y=683500
X861 4568 1 2 924 BUF1S $T=889080 618360 1 180 $X=886600 $Y=617980
X862 4780 1 2 4772 BUF1S $T=888460 648600 0 0 $X=888460 $Y=648220
X863 4762 1 2 4837 BUF1S $T=889080 709080 0 0 $X=889080 $Y=708700
X864 4169 1 2 940 BUF1S $T=890320 719160 1 0 $X=890320 $Y=713740
X865 897 1 2 4925 BUF1S $T=891560 588120 1 0 $X=891560 $Y=582700
X866 4820 1 2 4929 BUF1S $T=892180 588120 0 0 $X=892180 $Y=587740
X867 4733 1 2 4940 BUF1S $T=892180 709080 0 0 $X=892180 $Y=708700
X868 4883 1 2 4902 BUF1S $T=894040 668760 0 0 $X=894040 $Y=668380
X869 4799 1 2 4955 BUF1S $T=895900 628440 0 0 $X=895900 $Y=628060
X870 4822 1 2 4947 BUF1S $T=895900 638520 0 0 $X=895900 $Y=638140
X871 4672 1 2 4957 BUF1S $T=897140 658680 0 0 $X=897140 $Y=658300
X872 4744 1 2 4952 BUF1S $T=897140 678840 1 0 $X=897140 $Y=673420
X873 4888 1 2 4917 BUF1S $T=897760 567960 1 0 $X=897760 $Y=562540
X874 4951 1 2 4958 BUF1S $T=898380 688920 0 0 $X=898380 $Y=688540
X875 4760 1 2 4966 BUF1S $T=899000 628440 0 0 $X=899000 $Y=628060
X876 4954 1 2 4928 BUF1S $T=902720 547800 0 0 $X=902720 $Y=547420
X877 4660 1 2 4989 BUF1S $T=902720 658680 1 0 $X=902720 $Y=653260
X878 4935 1 2 962 BUF1S $T=904580 547800 1 0 $X=904580 $Y=542380
X879 4905 1 2 4976 BUF1S $T=904580 557880 0 0 $X=904580 $Y=557500
X880 4915 1 2 4990 BUF1S $T=905820 567960 1 0 $X=905820 $Y=562540
X881 4831 1 2 4959 BUF1S $T=906440 578040 1 0 $X=906440 $Y=572620
X882 5009 1 2 4936 BUF1S $T=908920 578040 0 0 $X=908920 $Y=577660
X883 4929 1 2 5039 BUF1S $T=910160 588120 0 0 $X=910160 $Y=587740
X884 4786 1 2 4998 BUF1S $T=915740 618360 0 180 $X=913260 $Y=612940
X885 4925 1 2 5037 BUF1S $T=915120 578040 1 0 $X=915120 $Y=572620
X886 968 1 2 4927 BUF1S $T=917600 699000 1 180 $X=915120 $Y=698620
X887 5058 1 2 4977 BUF1S $T=918840 578040 1 0 $X=918840 $Y=572620
X888 4870 1 2 4979 BUF1S $T=920080 699000 0 0 $X=920080 $Y=698620
X889 4912 1 2 5071 BUF1S $T=923180 557880 1 180 $X=920700 $Y=557500
X890 4870 1 2 5035 BUF1S $T=920700 699000 1 0 $X=920700 $Y=693580
X891 5008 1 2 5090 BUF1S $T=921320 567960 0 0 $X=921320 $Y=567580
X892 4943 1 2 5073 BUF1S $T=922560 578040 1 0 $X=922560 $Y=572620
X893 964 1 2 983 BUF1S $T=925040 719160 0 0 $X=925040 $Y=718780
X894 4979 1 2 5127 BUF1S $T=926280 719160 1 0 $X=926280 $Y=713740
X895 879 1 2 5151 BUF1S $T=931240 588120 0 0 $X=931240 $Y=587740
X896 4658 1 2 5149 BUF1S $T=934960 578040 1 0 $X=934960 $Y=572620
X897 5174 1 2 5186 BUF1S $T=936820 567960 0 0 $X=936820 $Y=567580
X898 4658 1 2 5207 BUF1S $T=941780 598200 1 0 $X=941780 $Y=592780
X899 5021 1 2 5217 BUF1S $T=941780 658680 1 0 $X=941780 $Y=653260
X900 5243 1 2 5082 BUF1S $T=947980 628440 0 180 $X=945500 $Y=623020
X901 5178 1 2 5275 BUF1S $T=949220 598200 1 0 $X=949220 $Y=592780
X902 5179 1 2 5260 BUF1S $T=951080 567960 0 0 $X=951080 $Y=567580
X903 5151 1 2 5194 BUF1S $T=951080 578040 1 0 $X=951080 $Y=572620
X904 975 1 2 5280 BUF1S $T=952320 699000 0 0 $X=952320 $Y=698620
X905 5288 1 2 5201 BUF1S $T=956660 578040 0 180 $X=954180 $Y=572620
X906 4877 1 2 5308 BUF1S $T=957900 578040 1 0 $X=957900 $Y=572620
X907 5127 1 2 5239 BUF1S $T=960380 709080 0 180 $X=957900 $Y=703660
X908 5282 1 2 5311 BUF1S $T=959760 567960 1 0 $X=959760 $Y=562540
X909 5288 1 2 1009 BUF1S $T=965960 567960 1 0 $X=965960 $Y=562540
X910 803 1 2 1020 BUF1S $T=966580 608280 0 0 $X=966580 $Y=607900
X911 5341 1 2 5288 BUF1S $T=970920 567960 0 180 $X=968440 $Y=562540
X912 5263 1 2 5313 BUF1S $T=969680 648600 1 0 $X=969680 $Y=643180
X913 5345 1 2 1028 BUF1S $T=970920 567960 1 0 $X=970920 $Y=562540
X914 1034 1 2 5312 BUF1S $T=980220 588120 0 180 $X=977740 $Y=582700
X915 5385 1 2 5374 BUF1S $T=980220 668760 0 180 $X=977740 $Y=663340
X916 5377 1 2 5348 BUF1S $T=977740 688920 0 0 $X=977740 $Y=688540
X917 5387 1 2 5400 BUF1S $T=980220 578040 1 0 $X=980220 $Y=572620
X918 5367 1 2 5371 BUF1S $T=983940 658680 0 0 $X=983940 $Y=658300
X919 5442 1 2 5414 BUF1S $T=988280 709080 1 0 $X=988280 $Y=703660
X920 5408 1 2 5448 BUF1S $T=991380 547800 1 180 $X=988900 $Y=547420
X921 5456 1 2 5341 BUF1S $T=991380 567960 1 180 $X=988900 $Y=567580
X922 1031 1 2 1061 BUF1S $T=990140 618360 0 0 $X=990140 $Y=617980
X923 5467 1 2 5407 BUF1S $T=993240 567960 0 180 $X=990760 $Y=562540
X924 5432 1 2 5478 BUF1S $T=991380 618360 1 0 $X=991380 $Y=612940
X925 1036 1 2 1068 BUF1S $T=991380 628440 0 0 $X=991380 $Y=628060
X926 1046 1 2 5477 BUF1S $T=991380 719160 1 0 $X=991380 $Y=713740
X927 5420 1 2 1072 BUF1S $T=993240 567960 1 0 $X=993240 $Y=562540
X928 5388 1 2 5449 BUF1S $T=993240 618360 0 0 $X=993240 $Y=617980
X929 5398 1 2 5346 BUF1S $T=995100 709080 1 0 $X=995100 $Y=703660
X930 5336 1 2 5383 BUF1S $T=998200 547800 0 0 $X=998200 $Y=547420
X931 5447 1 2 5492 BUF1S $T=1000680 709080 0 0 $X=1000680 $Y=708700
X932 5550 1 2 5450 BUF1S $T=1005020 688920 0 0 $X=1005020 $Y=688540
X933 5509 1 2 5525 BUF1S $T=1005640 618360 1 0 $X=1005640 $Y=612940
X934 5385 1 2 5579 BUF1S $T=1007500 668760 1 0 $X=1007500 $Y=663340
X935 5565 1 2 5577 BUF1S $T=1008120 567960 1 0 $X=1008120 $Y=562540
X936 5469 1 2 5578 BUF1S $T=1008120 678840 0 0 $X=1008120 $Y=678460
X937 5388 1 2 5584 BUF1S $T=1009360 628440 1 0 $X=1009360 $Y=623020
X938 5583 1 2 5598 BUF1S $T=1011220 567960 0 0 $X=1011220 $Y=567580
X939 5466 1 2 5612 BUF1S $T=1011220 648600 0 0 $X=1011220 $Y=648220
X940 5350 1 2 5608 BUF1S $T=1013080 638520 1 0 $X=1013080 $Y=633100
X941 5609 1 2 5354 BUF1S $T=1015560 678840 1 180 $X=1013080 $Y=678460
X942 5368 1 2 5610 BUF1S $T=1013080 699000 1 0 $X=1013080 $Y=693580
X943 5442 1 2 5605 BUF1S $T=1013080 709080 1 0 $X=1013080 $Y=703660
X944 5611 1 2 5474 BUF1S $T=1015560 709080 1 180 $X=1013080 $Y=708700
X945 5547 1 2 5597 BUF1S $T=1013700 567960 0 0 $X=1013700 $Y=567580
X946 5412 1 2 5625 BUF1S $T=1016180 628440 0 0 $X=1016180 $Y=628060
X947 5599 1 2 5629 BUF1S $T=1017420 598200 1 0 $X=1017420 $Y=592780
X948 5597 1 2 5638 BUF1S $T=1019900 578040 1 0 $X=1019900 $Y=572620
X949 5628 1 2 5648 BUF1S $T=1019900 709080 0 0 $X=1019900 $Y=708700
X950 5682 1 2 5554 BUF1S $T=1027960 699000 0 180 $X=1025480 $Y=693580
X951 5678 1 2 5686 BUF1S $T=1026100 699000 0 0 $X=1026100 $Y=698620
X952 5575 1 2 5702 BUF1S $T=1026720 588120 0 0 $X=1026720 $Y=587740
X953 5522 1 2 1109 BUF1S $T=1031680 588120 0 0 $X=1031680 $Y=587740
X954 5616 1 2 5609 BUF1S $T=1033540 688920 0 0 $X=1033540 $Y=688540
X955 5702 1 2 5683 BUF1S $T=1034160 598200 1 0 $X=1034160 $Y=592780
X956 5566 1 2 5717 BUF1S $T=1036020 578040 1 0 $X=1036020 $Y=572620
X957 5494 1 2 1110 BUF1S $T=1038500 588120 1 180 $X=1036020 $Y=587740
X958 5693 1 2 5672 BUF1S $T=1036640 668760 1 0 $X=1036640 $Y=663340
X959 5748 1 2 5421 BUF1S $T=1040360 648600 1 180 $X=1037880 $Y=648220
X960 5420 1 2 5751 BUF1S $T=1039740 588120 0 0 $X=1039740 $Y=587740
X961 5608 1 2 5771 BUF1S $T=1040980 638520 1 0 $X=1040980 $Y=633100
X962 5657 1 2 5724 BUF1S $T=1040980 709080 1 0 $X=1040980 $Y=703660
X963 1088 1 2 5744 BUF1S $T=1041600 567960 1 0 $X=1041600 $Y=562540
X964 5619 1 2 5763 BUF1S $T=1041600 567960 0 0 $X=1041600 $Y=567580
X965 5522 1 2 5782 BUF1S $T=1042840 588120 0 0 $X=1042840 $Y=587740
X966 5494 1 2 5774 BUF1S $T=1042840 608280 0 0 $X=1042840 $Y=607900
X967 5753 1 2 5770 BUF1S $T=1042840 678840 1 0 $X=1042840 $Y=673420
X968 5609 1 2 5748 BUF1S $T=1043460 678840 0 0 $X=1043460 $Y=678460
X969 5443 1 2 5794 BUF1S $T=1047180 557880 0 0 $X=1047180 $Y=557500
X970 5605 1 2 5806 BUF1S $T=1048420 699000 0 0 $X=1048420 $Y=698620
X971 5747 1 2 5616 BUF1S $T=1050900 709080 1 180 $X=1048420 $Y=708700
X972 5610 1 2 5813 BUF1S $T=1050280 709080 1 0 $X=1050280 $Y=703660
X973 5702 1 2 5822 BUF1S $T=1051520 578040 1 0 $X=1051520 $Y=572620
X974 5625 1 2 5838 BUF1S $T=1052140 618360 0 0 $X=1052140 $Y=617980
X975 5747 1 2 1107 BUF1S $T=1055860 709080 0 180 $X=1053380 $Y=703660
X976 5612 1 2 5845 BUF1S $T=1055240 658680 1 0 $X=1055240 $Y=653260
X977 5448 1 2 5842 BUF1S $T=1055860 537720 0 0 $X=1055860 $Y=537340
X978 5747 1 2 5865 BUF1S $T=1057100 709080 0 0 $X=1057100 $Y=708700
X979 5863 1 2 5765 BUF1S $T=1061440 618360 1 180 $X=1058960 $Y=617980
X980 5857 1 2 5863 BUF1S $T=1058960 658680 1 0 $X=1058960 $Y=653260
X981 5858 1 2 5732 BUF1S $T=1059580 678840 1 0 $X=1059580 $Y=673420
X982 5757 1 2 5818 BUF1S $T=1059580 688920 0 0 $X=1059580 $Y=688540
X983 5754 1 2 5906 BUF1S $T=1070740 678840 1 0 $X=1070740 $Y=673420
X984 5879 1 2 5869 BUF1S $T=1071980 658680 1 0 $X=1071980 $Y=653260
X985 5886 1 2 5914 BUF1S $T=1073840 618360 1 0 $X=1073840 $Y=612940
X986 5974 1 2 5991 BUF1S $T=1084380 628440 1 0 $X=1084380 $Y=623020
X987 5937 1 2 1143 BUF1S $T=1088720 547800 1 0 $X=1088720 $Y=542380
X988 5936 1 2 5989 BUF1S $T=1091820 709080 0 180 $X=1089340 $Y=703660
X989 5990 1 2 6054 BUF1S $T=1095540 598200 1 0 $X=1095540 $Y=592780
X990 6001 1 2 5975 BUF1S $T=1098020 668760 0 0 $X=1098020 $Y=668380
X991 6071 1 2 6094 BUF1S $T=1101120 688920 0 0 $X=1101120 $Y=688540
X992 5936 1 2 1175 BUF1S $T=1105460 709080 0 0 $X=1105460 $Y=708700
X993 5995 1 2 6138 BUF1S $T=1109180 608280 0 0 $X=1109180 $Y=607900
X994 6139 1 2 6164 BUF1S $T=1112900 668760 0 0 $X=1112900 $Y=668380
X995 1146 1 2 1183 BUF1S $T=1116620 719160 1 0 $X=1116620 $Y=713740
X996 6159 1 2 1179 BUF1S $T=1123440 537720 0 0 $X=1123440 $Y=537340
X997 6178 1 2 6131 BUF1S $T=1129020 648600 1 180 $X=1126540 $Y=648220
X998 1175 1 2 6178 BUF1S $T=1126540 699000 0 0 $X=1126540 $Y=698620
X999 1238 1 2 1253 DELB $T=221960 709080 0 0 $X=221960 $Y=708700
X1000 1338 1 2 1332 DELB $T=236840 688920 1 0 $X=236840 $Y=683500
X1001 1339 1 2 18 DELB $T=238700 709080 0 0 $X=238700 $Y=708700
X1002 1507 1 2 1529 DELB $T=267840 567960 0 0 $X=267840 $Y=567580
X1003 1841 1 2 1894 DELB $T=347200 678840 1 0 $X=347200 $Y=673420
X1004 2104 1 2 2115 DELB $T=387500 598200 1 0 $X=387500 $Y=592780
X1005 2195 1 2 2233 DELB $T=405480 628440 1 0 $X=405480 $Y=623020
X1006 2312 1 2 2239 DELB $T=419120 598200 1 0 $X=419120 $Y=592780
X1007 2313 1 2 2347 DELB $T=422220 628440 0 0 $X=422220 $Y=628060
X1008 2358 1 2 2360 DELB $T=426560 598200 1 0 $X=426560 $Y=592780
X1009 288 1 2 293 DELB $T=473060 719160 0 0 $X=473060 $Y=718780
X1010 2697 1 2 2711 DELB $T=484220 688920 0 0 $X=484220 $Y=688540
X1011 2721 1 2 2756 DELB $T=489800 709080 0 0 $X=489800 $Y=708700
X1012 328 1 2 337 DELB $T=499720 537720 0 0 $X=499720 $Y=537340
X1013 2811 1 2 2864 DELB $T=513980 699000 0 0 $X=513980 $Y=698620
X1014 2869 1 2 2901 DELB $T=515840 648600 1 0 $X=515840 $Y=643180
X1015 2883 1 2 2912 DELB $T=516460 658680 0 0 $X=516460 $Y=658300
X1016 370 1 2 376 DELB $T=522040 678840 0 0 $X=522040 $Y=678460
X1017 2942 1 2 2958 DELB $T=530100 547800 0 0 $X=530100 $Y=547420
X1018 2976 1 2 3005 DELB $T=533200 638520 1 0 $X=533200 $Y=633100
X1019 392 1 2 400 DELB $T=536920 688920 0 0 $X=536920 $Y=688540
X1020 2965 1 2 3011 DELB $T=538160 709080 1 0 $X=538160 $Y=703660
X1021 3019 1 2 3014 DELB $T=539400 547800 0 0 $X=539400 $Y=547420
X1022 2984 1 2 3029 DELB $T=540640 719160 0 0 $X=540640 $Y=718780
X1023 409 1 2 3075 DELB $T=547460 709080 1 0 $X=547460 $Y=703660
X1024 3016 1 2 3087 DELB $T=551800 699000 0 0 $X=551800 $Y=698620
X1025 3102 1 2 3117 DELB $T=555520 668760 1 0 $X=555520 $Y=663340
X1026 3093 1 2 3109 DELB $T=557380 699000 0 0 $X=557380 $Y=698620
X1027 3121 1 2 3146 DELB $T=561100 628440 1 0 $X=561100 $Y=623020
X1028 3059 1 2 3086 DELB $T=565440 699000 1 0 $X=565440 $Y=693580
X1029 453 1 2 465 DELB $T=567920 668760 0 0 $X=567920 $Y=668380
X1030 464 1 2 476 DELB $T=572260 658680 1 0 $X=572260 $Y=653260
X1031 3175 1 2 3205 DELB $T=572880 588120 1 0 $X=572880 $Y=582700
X1032 472 1 2 487 DELB $T=577840 699000 1 0 $X=577840 $Y=693580
X1033 490 1 2 498 DELB $T=583420 648600 0 0 $X=583420 $Y=648220
X1034 3259 1 2 3282 DELB $T=587760 608280 1 0 $X=587760 $Y=602860
X1035 3293 1 2 3312 DELB $T=593960 588120 1 0 $X=593960 $Y=582700
X1036 513 1 2 523 DELB $T=594580 608280 0 0 $X=594580 $Y=607900
X1037 3378 1 2 3399 DELB $T=610700 618360 1 0 $X=610700 $Y=612940
X1038 3389 1 2 3416 DELB $T=613800 578040 0 0 $X=613800 $Y=577660
X1039 583 1 2 590 DELB $T=618760 699000 0 0 $X=618760 $Y=698620
X1040 3343 1 2 3427 DELB $T=619380 688920 1 0 $X=619380 $Y=683500
X1041 3476 1 2 3506 DELB $T=629300 557880 1 0 $X=629300 $Y=552460
X1042 3496 1 2 3529 DELB $T=631780 567960 1 0 $X=631780 $Y=562540
X1043 3557 1 2 3545 DELB $T=644180 588120 1 0 $X=644180 $Y=582700
X1044 3558 1 2 3593 DELB $T=647280 648600 1 0 $X=647280 $Y=643180
X1045 640 1 2 644 DELB $T=649140 719160 0 0 $X=649140 $Y=718780
X1046 3586 1 2 3612 DELB $T=652240 678840 1 0 $X=652240 $Y=673420
X1047 3614 1 2 3642 DELB $T=657820 608280 0 0 $X=657820 $Y=607900
X1048 3643 1 2 3683 DELB $T=657820 658680 0 0 $X=657820 $Y=658300
X1049 3631 1 2 3661 DELB $T=658440 658680 1 0 $X=658440 $Y=653260
X1050 3662 1 2 3621 DELB $T=660920 688920 1 0 $X=660920 $Y=683500
X1051 3691 1 2 3690 DELB $T=664640 547800 0 0 $X=664640 $Y=547420
X1052 642 1 2 3641 DELB $T=666500 709080 1 0 $X=666500 $Y=703660
X1053 3703 1 2 3699 DELB $T=667120 608280 0 0 $X=667120 $Y=607900
X1054 3710 1 2 3733 DELB $T=668360 567960 0 0 $X=668360 $Y=567580
X1055 3719 1 2 3720 DELB $T=669600 688920 1 0 $X=669600 $Y=683500
X1056 3779 1 2 3799 DELB $T=680760 678840 0 0 $X=680760 $Y=678460
X1057 3780 1 2 3772 DELB $T=681380 578040 1 0 $X=681380 $Y=572620
X1058 3773 1 2 3781 DELB $T=683860 608280 0 0 $X=683860 $Y=607900
X1059 3793 1 2 3814 DELB $T=684480 638520 1 0 $X=684480 $Y=633100
X1060 3805 1 2 3807 DELB $T=686340 699000 1 0 $X=686340 $Y=693580
X1061 3796 1 2 3783 DELB $T=686960 668760 0 0 $X=686960 $Y=668380
X1062 3787 1 2 3836 DELB $T=688200 578040 1 0 $X=688200 $Y=572620
X1063 3827 1 2 3823 DELB $T=693160 648600 1 0 $X=693160 $Y=643180
X1064 3850 1 2 3872 DELB $T=698740 618360 1 0 $X=698740 $Y=612940
X1065 3815 1 2 3863 DELB $T=699980 658680 0 0 $X=699980 $Y=658300
X1066 3898 1 2 3901 DELB $T=704940 668760 1 0 $X=704940 $Y=663340
X1067 3945 1 2 3964 DELB $T=715480 557880 1 0 $X=715480 $Y=552460
X1068 3963 1 2 3965 DELB $T=719200 688920 0 0 $X=719200 $Y=688540
X1069 3969 1 2 3962 DELB $T=720440 688920 1 0 $X=720440 $Y=683500
X1070 3976 1 2 3975 DELB $T=721680 578040 0 0 $X=721680 $Y=577660
X1071 3990 1 2 4014 DELB $T=724160 648600 0 0 $X=724160 $Y=648220
X1072 4003 1 2 4028 DELB $T=729120 608280 0 0 $X=729120 $Y=607900
X1073 3993 1 2 3989 DELB $T=730980 638520 0 0 $X=730980 $Y=638140
X1074 3973 1 2 4016 DELB $T=739040 608280 1 0 $X=739040 $Y=602860
X1075 4063 1 2 4074 DELB $T=743380 588120 1 0 $X=743380 $Y=582700
X1076 4086 1 2 4118 DELB $T=743380 699000 0 0 $X=743380 $Y=698620
X1077 4001 1 2 4078 DELB $T=744620 678840 0 0 $X=744620 $Y=678460
X1078 768 1 2 773 DELB $T=748340 547800 1 0 $X=748340 $Y=542380
X1079 4127 1 2 4150 DELB $T=750820 709080 0 0 $X=750820 $Y=708700
X1080 4128 1 2 4131 DELB $T=751440 618360 0 0 $X=751440 $Y=617980
X1081 4130 1 2 4159 DELB $T=752060 678840 0 0 $X=752060 $Y=678460
X1082 4137 1 2 4132 DELB $T=756400 628440 1 0 $X=756400 $Y=623020
X1083 4160 1 2 4155 DELB $T=757020 688920 0 0 $X=757020 $Y=688540
X1084 4158 1 2 4149 DELB $T=761360 678840 1 0 $X=761360 $Y=673420
X1085 4193 1 2 4192 DELB $T=761980 648600 1 0 $X=761980 $Y=643180
X1086 4199 1 2 4198 DELB $T=763220 688920 0 0 $X=763220 $Y=688540
X1087 4142 1 2 4196 DELB $T=766320 547800 1 0 $X=766320 $Y=542380
X1088 4227 1 2 4228 DELB $T=769420 648600 1 0 $X=769420 $Y=643180
X1089 4136 1 2 4181 DELB $T=773760 658680 0 0 $X=773760 $Y=658300
X1090 4270 1 2 4249 DELB $T=778100 567960 1 0 $X=778100 $Y=562540
X1091 4256 1 2 4271 DELB $T=778100 678840 0 0 $X=778100 $Y=678460
X1092 4274 1 2 4273 DELB $T=778720 628440 1 0 $X=778720 $Y=623020
X1093 4301 1 2 4310 DELB $T=784920 678840 0 0 $X=784920 $Y=678460
X1094 4300 1 2 4335 DELB $T=789880 668760 1 0 $X=789880 $Y=663340
X1095 4257 1 2 4246 DELB $T=790500 547800 1 0 $X=790500 $Y=542380
X1096 4284 1 2 4318 DELB $T=792360 699000 0 0 $X=792360 $Y=698620
X1097 4344 1 2 4380 DELB $T=794220 628440 0 0 $X=794220 $Y=628060
X1098 4339 1 2 4345 DELB $T=796080 598200 0 0 $X=796080 $Y=597820
X1099 4351 1 2 4370 DELB $T=797940 598200 1 0 $X=797940 $Y=592780
X1100 4373 1 2 4409 DELB $T=804760 668760 0 0 $X=804760 $Y=668380
X1101 4355 1 2 4401 DELB $T=806620 588120 0 0 $X=806620 $Y=587740
X1102 4376 1 2 4435 DELB $T=813440 547800 0 0 $X=813440 $Y=547420
X1103 4383 1 2 4410 DELB $T=815300 678840 0 0 $X=815300 $Y=678460
X1104 4361 1 2 4358 DELB $T=817160 638520 1 0 $X=817160 $Y=633100
X1105 4337 1 2 4439 DELB $T=818400 588120 1 0 $X=818400 $Y=582700
X1106 4520 1 2 4555 DELB $T=825840 658680 0 0 $X=825840 $Y=658300
X1107 4512 1 2 4548 DELB $T=827080 588120 1 0 $X=827080 $Y=582700
X1108 4535 1 2 4567 DELB $T=828320 688920 1 0 $X=828320 $Y=683500
X1109 4559 1 2 4553 DELB $T=830800 557880 1 0 $X=830800 $Y=552460
X1110 4572 1 2 4580 DELB $T=835140 668760 0 0 $X=835140 $Y=668380
X1111 4569 1 2 4574 DELB $T=837000 588120 1 0 $X=837000 $Y=582700
X1112 4560 1 2 4554 DELB $T=837000 638520 1 0 $X=837000 $Y=633100
X1113 4334 1 2 4377 DELB $T=837620 547800 1 0 $X=837620 $Y=542380
X1114 4536 1 2 4571 DELB $T=841960 578040 0 0 $X=841960 $Y=577660
X1115 4624 1 2 4623 DELB $T=841960 678840 0 0 $X=841960 $Y=678460
X1116 4575 1 2 4565 DELB $T=842580 608280 1 0 $X=842580 $Y=602860
X1117 883 1 2 888 DELB $T=843200 547800 1 0 $X=843200 $Y=542380
X1118 4606 1 2 4622 DELB $T=845060 618360 0 0 $X=845060 $Y=617980
X1119 4613 1 2 4636 DELB $T=846300 588120 1 0 $X=846300 $Y=582700
X1120 4549 1 2 4576 DELB $T=856220 658680 1 0 $X=856220 $Y=653260
X1121 4693 1 2 4717 DELB $T=858080 688920 1 0 $X=858080 $Y=683500
X1122 4724 1 2 4702 DELB $T=861800 608280 1 0 $X=861800 $Y=602860
X1123 908 1 2 4773 DELB $T=863040 719160 0 0 $X=863040 $Y=718780
X1124 4734 1 2 4756 DELB $T=865520 578040 0 0 $X=865520 $Y=577660
X1125 4774 1 2 4776 DELB $T=868000 608280 1 0 $X=868000 $Y=602860
X1126 4782 1 2 4796 DELB $T=869240 648600 1 0 $X=869240 $Y=643180
X1127 4791 1 2 4812 DELB $T=874820 668760 0 0 $X=874820 $Y=668380
X1128 4842 1 2 4879 DELB $T=880400 668760 0 0 $X=880400 $Y=668380
X1129 4808 1 2 4811 DELB $T=882260 598200 1 0 $X=882260 $Y=592780
X1130 4518 1 2 4603 DELB $T=887220 557880 1 0 $X=887220 $Y=552460
X1131 4899 1 2 4865 DELB $T=891560 608280 0 0 $X=891560 $Y=607900
X1132 942 1 2 4946 DELB $T=896520 678840 0 0 $X=896520 $Y=678460
X1133 946 1 2 956 DELB $T=899000 688920 1 0 $X=899000 $Y=683500
X1134 4956 1 2 4960 DELB $T=899620 608280 0 0 $X=899620 $Y=607900
X1135 4800 1 2 4854 DELB $T=903340 567960 0 0 $X=903340 $Y=567580
X1136 959 1 2 5022 DELB $T=905200 537720 0 0 $X=905200 $Y=537340
X1137 4920 1 2 4993 DELB $T=905820 608280 0 0 $X=905820 $Y=607900
X1138 4987 1 2 4978 DELB $T=907060 628440 0 0 $X=907060 $Y=628060
X1139 5038 1 2 5062 DELB $T=912640 578040 0 0 $X=912640 $Y=577660
X1140 5015 1 2 5051 DELB $T=914500 628440 0 0 $X=914500 $Y=628060
X1141 4953 1 2 4995 DELB $T=915740 608280 0 0 $X=915740 $Y=607900
X1142 5060 1 2 5081 DELB $T=916360 588120 1 0 $X=916360 $Y=582700
X1143 5068 1 2 5042 DELB $T=920700 618360 1 0 $X=920700 $Y=612940
X1144 5017 1 2 5061 DELB $T=920700 688920 1 0 $X=920700 $Y=683500
X1145 5107 1 2 5130 DELB $T=925040 578040 1 0 $X=925040 $Y=572620
X1146 5125 1 2 5115 DELB $T=927520 678840 1 0 $X=927520 $Y=673420
X1147 5087 1 2 5096 DELB $T=932480 638520 1 0 $X=932480 $Y=633100
X1148 5148 1 2 5162 DELB $T=934340 557880 1 0 $X=934340 $Y=552460
X1149 5173 1 2 5209 DELB $T=939300 567960 0 0 $X=939300 $Y=567580
X1150 5132 1 2 5181 DELB $T=939300 688920 1 0 $X=939300 $Y=683500
X1151 5168 1 2 5198 DELB $T=939920 638520 0 0 $X=939920 $Y=638140
X1152 5182 1 2 5200 DELB $T=945500 567960 1 0 $X=945500 $Y=562540
X1153 5251 1 2 5296 DELB $T=952940 588120 1 0 $X=952940 $Y=582700
X1154 5270 1 2 5297 DELB $T=953560 557880 0 0 $X=953560 $Y=557500
X1155 5237 1 2 5262 DELB $T=954800 678840 1 0 $X=954800 $Y=673420
X1156 5302 1 2 5320 DELB $T=969060 608280 0 0 $X=969060 $Y=607900
X1157 5342 1 2 5361 DELB $T=970300 598200 0 0 $X=970300 $Y=597820
X1158 4677 1 2 4707 DELB $T=973400 578040 1 0 $X=973400 $Y=572620
X1159 5293 1 2 5365 DELB $T=974020 588120 0 0 $X=974020 $Y=587740
X1160 5391 1 2 5394 DELB $T=980220 688920 0 0 $X=980220 $Y=688540
X1161 5010 1 2 5063 DELB $T=982080 678840 1 0 $X=982080 $Y=673420
X1162 5384 1 2 5416 DELB $T=984560 628440 1 0 $X=984560 $Y=623020
X1163 1041 1 2 1054 DELB $T=985180 537720 0 0 $X=985180 $Y=537340
X1164 1043 1 2 1057 DELB $T=985180 699000 0 0 $X=985180 $Y=698620
X1165 5397 1 2 5390 DELB $T=987040 668760 0 0 $X=987040 $Y=668380
X1166 5409 1 2 5389 DELB $T=988900 658680 0 0 $X=988900 $Y=658300
X1167 5462 1 2 5461 DELB $T=991380 699000 0 0 $X=991380 $Y=698620
X1168 5476 1 2 5485 DELB $T=995100 578040 0 0 $X=995100 $Y=577660
X1169 5472 1 2 5503 DELB $T=996960 699000 0 0 $X=996960 $Y=698620
X1170 5500 1 2 5535 DELB $T=998820 658680 1 0 $X=998820 $Y=653260
X1171 5431 1 2 5465 DELB $T=998820 668760 1 0 $X=998820 $Y=663340
X1172 5533 1 2 5532 DELB $T=1003160 699000 0 0 $X=1003160 $Y=698620
X1173 4670 1 2 4715 DELB $T=1005020 658680 0 0 $X=1005020 $Y=658300
X1174 5558 1 2 5559 DELB $T=1006880 588120 1 0 $X=1006880 $Y=582700
X1175 5562 1 2 5557 DELB $T=1007500 709080 0 0 $X=1007500 $Y=708700
X1176 5570 1 2 5569 DELB $T=1008740 618360 1 0 $X=1008740 $Y=612940
X1177 5585 1 2 5620 DELB $T=1011220 658680 0 0 $X=1011220 $Y=658300
X1178 5588 1 2 5603 DELB $T=1014320 557880 0 0 $X=1014320 $Y=557500
X1179 5602 1 2 5647 DELB $T=1021140 688920 0 0 $X=1021140 $Y=688540
X1180 5592 1 2 5622 DELB $T=1022380 567960 1 0 $X=1022380 $Y=562540
X1181 5655 1 2 5630 DELB $T=1023620 638520 1 0 $X=1023620 $Y=633100
X1182 5698 1 2 5658 DELB $T=1029820 618360 0 0 $X=1029820 $Y=617980
X1183 5688 1 2 5699 DELB $T=1029820 709080 1 0 $X=1029820 $Y=703660
X1184 5689 1 2 5703 DELB $T=1030440 578040 0 0 $X=1030440 $Y=577660
X1185 5700 1 2 5651 DELB $T=1036640 628440 1 0 $X=1036640 $Y=623020
X1186 5736 1 2 5767 DELB $T=1043460 709080 1 0 $X=1043460 $Y=703660
X1187 5738 1 2 5752 DELB $T=1047180 618360 1 0 $X=1047180 $Y=612940
X1188 5766 1 2 5789 DELB $T=1049660 638520 0 0 $X=1049660 $Y=638140
X1189 5756 1 2 5776 DELB $T=1049660 658680 1 0 $X=1049660 $Y=653260
X1190 1122 1 2 5835 DELB $T=1050900 709080 0 0 $X=1050900 $Y=708700
X1191 5823 1 2 5852 DELB $T=1054620 668760 0 0 $X=1054620 $Y=668380
X1192 5833 1 2 5832 DELB $T=1054620 699000 0 0 $X=1054620 $Y=698620
X1193 1124 1 2 5793 DELB $T=1058340 537720 0 0 $X=1058340 $Y=537340
X1194 5846 1 2 5875 DELB $T=1058340 557880 0 0 $X=1058340 $Y=557500
X1195 5811 1 2 5860 DELB $T=1058960 638520 0 0 $X=1058960 $Y=638140
X1196 5872 1 2 5898 DELB $T=1062680 658680 1 0 $X=1062680 $Y=653260
X1197 5824 1 2 5850 DELB $T=1063300 547800 1 0 $X=1063300 $Y=542380
X1198 5837 1 2 5873 DELB $T=1063300 668760 0 0 $X=1063300 $Y=668380
X1199 5884 1 2 5900 DELB $T=1065780 578040 1 0 $X=1065780 $Y=572620
X1200 5848 1 2 5896 DELB $T=1067640 638520 0 0 $X=1067640 $Y=638140
X1201 5908 1 2 5931 DELB $T=1069500 547800 1 0 $X=1069500 $Y=542380
X1202 5909 1 2 5912 DELB $T=1069500 699000 1 0 $X=1069500 $Y=693580
X1203 5856 1 2 5862 DELB $T=1071360 608280 0 0 $X=1071360 $Y=607900
X1204 5938 1 2 5959 DELB $T=1075700 688920 0 0 $X=1075700 $Y=688540
X1205 1141 1 2 1159 DELB $T=1082520 719160 0 0 $X=1082520 $Y=718780
X1206 5978 1 2 5965 DELB $T=1084380 709080 1 0 $X=1084380 $Y=703660
X1207 1161 1 2 1167 DELB $T=1091820 719160 0 0 $X=1091820 $Y=718780
X1208 6000 1 2 5980 DELB $T=1098020 628440 0 0 $X=1098020 $Y=628060
X1209 6037 1 2 6065 DELB $T=1099880 598200 1 0 $X=1099880 $Y=592780
X1210 6070 1 2 6090 DELB $T=1103600 567960 1 0 $X=1103600 $Y=562540
X1211 6103 1 2 6127 DELB $T=1106080 598200 1 0 $X=1106080 $Y=592780
X1212 6091 1 2 6136 DELB $T=1119720 588120 1 0 $X=1119720 $Y=582700
X1213 6113 1 2 6179 DELB $T=1121580 547800 0 0 $X=1121580 $Y=547420
X1214 6129 1 2 6174 DELB $T=1122200 658680 1 0 $X=1122200 $Y=653260
X1215 1188 1 2 1191 DELB $T=1124680 709080 0 0 $X=1124680 $Y=708700
X1216 1254 1 2 1279 DELA $T=221960 567960 0 0 $X=221960 $Y=567580
X1217 1263 1 2 1245 DELA $T=224440 557880 1 0 $X=224440 $Y=552460
X1218 1276 1 2 1298 DELA $T=226300 598200 0 0 $X=226300 $Y=597820
X1219 1240 1 2 1283 DELA $T=234980 628440 1 0 $X=234980 $Y=623020
X1220 1327 1 2 1328 DELA $T=235600 557880 0 0 $X=235600 $Y=557500
X1221 1372 1 2 1417 DELA $T=245520 709080 0 0 $X=245520 $Y=708700
X1222 1434 1 2 1461 DELA $T=253580 567960 1 0 $X=253580 $Y=562540
X1223 1427 1 2 50 DELA $T=254820 547800 0 0 $X=254820 $Y=547420
X1224 1514 1 2 1515 DELA $T=269080 628440 0 0 $X=269080 $Y=628060
X1225 1510 1 2 1519 DELA $T=271560 598200 0 0 $X=271560 $Y=597820
X1226 1533 1 2 1554 DELA $T=275900 648600 1 0 $X=275900 $Y=643180
X1227 1582 1 2 1588 DELA $T=282100 578040 0 0 $X=282100 $Y=577660
X1228 1591 1 2 1596 DELA $T=283340 648600 1 0 $X=283340 $Y=643180
X1229 1606 1 2 1627 DELA $T=285820 588120 0 0 $X=285820 $Y=587740
X1230 1539 1 2 1613 DELA $T=286440 547800 0 0 $X=286440 $Y=547420
X1231 1617 1 2 1602 DELA $T=288300 578040 0 0 $X=288300 $Y=577660
X1232 1584 1 2 1561 DELA $T=288920 618360 1 0 $X=288920 $Y=612940
X1233 1697 1 2 1722 DELA $T=305660 709080 0 0 $X=305660 $Y=708700
X1234 1707 1 2 1700 DELA $T=306280 628440 0 0 $X=306280 $Y=628060
X1235 1654 1 2 1698 DELA $T=308140 578040 0 0 $X=308140 $Y=577660
X1236 1739 1 2 1767 DELA $T=311240 638520 0 0 $X=311240 $Y=638140
X1237 123 1 2 1756 DELA $T=313720 709080 1 0 $X=313720 $Y=703660
X1238 1765 1 2 1764 DELA $T=315580 578040 0 0 $X=315580 $Y=577660
X1239 1782 1 2 1777 DELA $T=318060 628440 0 0 $X=318060 $Y=628060
X1240 1759 1 2 1750 DELA $T=318680 588120 1 0 $X=318680 $Y=582700
X1241 132 1 2 1789 DELA $T=319300 709080 0 0 $X=319300 $Y=708700
X1242 1815 1 2 1837 DELA $T=324880 628440 0 0 $X=324880 $Y=628060
X1243 1826 1 2 1827 DELA $T=326740 648600 1 0 $X=326740 $Y=643180
X1244 1810 1 2 1828 DELA $T=326740 688920 1 0 $X=326740 $Y=683500
X1245 1847 1 2 1875 DELA $T=332320 658680 1 0 $X=332320 $Y=653260
X1246 1880 1 2 1879 DELA $T=339760 598200 1 0 $X=339760 $Y=592780
X1247 1881 1 2 1902 DELA $T=339760 648600 0 0 $X=339760 $Y=648220
X1248 1887 1 2 1918 DELA $T=341000 618360 0 0 $X=341000 $Y=617980
X1249 1927 1 2 1953 DELA $T=347820 598200 1 0 $X=347820 $Y=592780
X1250 1934 1 2 1933 DELA $T=348440 658680 0 0 $X=348440 $Y=658300
X1251 1946 1 2 1915 DELA $T=352160 628440 0 0 $X=352160 $Y=628060
X1252 1956 1 2 1959 DELA $T=353400 598200 0 0 $X=353400 $Y=597820
X1253 1991 1 2 2017 DELA $T=361460 628440 0 0 $X=361460 $Y=628060
X1254 1996 1 2 2025 DELA $T=363320 598200 1 0 $X=363320 $Y=592780
X1255 1869 1 2 1998 DELA $T=363320 658680 0 0 $X=363320 $Y=658300
X1256 2016 1 2 2036 DELA $T=366420 618360 1 0 $X=366420 $Y=612940
X1257 2018 1 2 2050 DELA $T=370760 638520 0 0 $X=370760 $Y=638140
X1258 2045 1 2 2055 DELA $T=380060 658680 1 0 $X=380060 $Y=653260
X1259 2057 1 2 2087 DELA $T=385020 567960 1 0 $X=385020 $Y=562540
X1260 2126 1 2 2140 DELA $T=386880 658680 1 0 $X=386880 $Y=653260
X1261 2153 1 2 2147 DELA $T=391840 578040 0 0 $X=391840 $Y=577660
X1262 2167 1 2 2191 DELA $T=393080 598200 1 0 $X=393080 $Y=592780
X1263 2131 1 2 2119 DELA $T=393080 628440 0 0 $X=393080 $Y=628060
X1264 2158 1 2 2185 DELA $T=393080 658680 0 0 $X=393080 $Y=658300
X1265 2171 1 2 2193 DELA $T=393700 618360 0 0 $X=393700 $Y=617980
X1266 2179 1 2 2156 DELA $T=395560 608280 1 0 $X=395560 $Y=602860
X1267 2202 1 2 2229 DELA $T=399280 628440 0 0 $X=399280 $Y=628060
X1268 2194 1 2 2182 DELA $T=400520 648600 1 0 $X=400520 $Y=643180
X1269 2215 1 2 2251 DELA $T=406100 598200 1 0 $X=406100 $Y=592780
X1270 2282 1 2 2304 DELA $T=414160 598200 1 0 $X=414160 $Y=592780
X1271 2257 1 2 2283 DELA $T=414160 618360 1 0 $X=414160 $Y=612940
X1272 2272 1 2 2309 DELA $T=416640 658680 0 0 $X=416640 $Y=658300
X1273 2292 1 2 2328 DELA $T=417260 628440 0 0 $X=417260 $Y=628060
X1274 2363 1 2 2341 DELA $T=427800 567960 0 0 $X=427800 $Y=567580
X1275 2390 1 2 2399 DELA $T=435860 598200 1 0 $X=435860 $Y=592780
X1276 238 1 2 2424 DELA $T=448880 557880 0 0 $X=448880 $Y=557500
X1277 2497 1 2 2461 DELA $T=449500 588120 1 0 $X=449500 $Y=582700
X1278 284 1 2 287 DELA $T=468100 719160 0 0 $X=468100 $Y=718780
X1279 310 1 2 318 DELA $T=486080 709080 1 0 $X=486080 $Y=703660
X1280 2830 1 2 2856 DELA $T=507780 668760 0 0 $X=507780 $Y=668380
X1281 2851 1 2 2877 DELA $T=511500 658680 0 0 $X=511500 $Y=658300
X1282 2931 1 2 2955 DELA $T=524520 678840 1 0 $X=524520 $Y=673420
X1283 414 1 2 421 DELA $T=549320 628440 1 0 $X=549320 $Y=623020
X1284 416 1 2 428 DELA $T=552420 648600 0 0 $X=552420 $Y=648220
X1285 417 1 2 430 DELA $T=553660 678840 0 0 $X=553660 $Y=678460
X1286 424 1 2 435 DELA $T=555520 618360 0 0 $X=555520 $Y=617980
X1287 440 1 2 451 DELA $T=562960 668760 0 0 $X=562960 $Y=668380
X1288 450 1 2 463 DELA $T=567300 648600 0 0 $X=567300 $Y=648220
X1289 3178 1 2 3183 DELA $T=572880 699000 1 0 $X=572880 $Y=693580
X1290 3194 1 2 3214 DELA $T=575360 608280 1 0 $X=575360 $Y=602860
X1291 3208 1 2 3222 DELA $T=577840 628440 1 0 $X=577840 $Y=623020
X1292 480 1 2 489 DELA $T=578460 648600 0 0 $X=578460 $Y=648220
X1293 485 1 2 494 DELA $T=582180 567960 0 0 $X=582180 $Y=567580
X1294 3266 1 2 3290 DELA $T=588380 588120 0 0 $X=588380 $Y=587740
X1295 500 1 2 509 DELA $T=589000 658680 1 0 $X=589000 $Y=653260
X1296 507 1 2 519 DELA $T=591480 628440 0 0 $X=591480 $Y=628060
X1297 3281 1 2 3299 DELA $T=592100 578040 1 0 $X=592100 $Y=572620
X1298 3294 1 2 3309 DELA $T=593960 608280 1 0 $X=593960 $Y=602860
X1299 515 1 2 525 DELA $T=594580 699000 1 0 $X=594580 $Y=693580
X1300 520 1 2 532 DELA $T=596440 598200 1 0 $X=596440 $Y=592780
X1301 528 1 2 541 DELA $T=599540 678840 1 0 $X=599540 $Y=673420
X1302 3336 1 2 3359 DELA $T=603260 567960 0 0 $X=603260 $Y=567580
X1303 3344 1 2 3372 DELA $T=605120 588120 1 0 $X=605120 $Y=582700
X1304 556 1 2 567 DELA $T=608840 678840 1 0 $X=608840 $Y=673420
X1305 564 1 2 578 DELA $T=611940 638520 0 0 $X=611940 $Y=638140
X1306 570 1 2 581 DELA $T=614420 598200 0 0 $X=614420 $Y=597820
X1307 3449 1 2 3477 DELA $T=624960 578040 1 0 $X=624960 $Y=572620
X1308 3461 1 2 3491 DELA $T=626820 567960 1 0 $X=626820 $Y=562540
X1309 625 1 2 634 DELA $T=639840 648600 0 0 $X=639840 $Y=648220
X1310 3599 1 2 3623 DELA $T=649760 598200 1 0 $X=649760 $Y=592780
X1311 3611 1 2 3635 DELA $T=651620 638520 0 0 $X=651620 $Y=638140
X1312 3625 1 2 3655 DELA $T=654100 628440 1 0 $X=654100 $Y=623020
X1313 3653 1 2 3685 DELA $T=659680 547800 0 0 $X=659680 $Y=547420
X1314 3696 1 2 3704 DELA $T=667120 658680 1 0 $X=667120 $Y=653260
X1315 3762 1 2 3775 DELA $T=677660 567960 0 0 $X=677660 $Y=567580
X1316 3881 1 2 3867 DELA $T=703700 547800 1 0 $X=703700 $Y=542380
X1317 3907 1 2 3911 DELA $T=719200 628440 0 0 $X=719200 $Y=628060
X1318 765 1 2 769 DELA $T=745860 709080 0 0 $X=745860 $Y=708700
X1319 4234 1 2 4266 DELA $T=779960 699000 1 0 $X=779960 $Y=693580
X1320 4491 1 2 4511 DELA $T=820880 709080 0 0 $X=820880 $Y=708700
X1321 4656 1 2 4626 DELA $T=848160 678840 0 0 $X=848160 $Y=678460
X1322 4686 1 2 4665 DELA $T=855600 668760 1 0 $X=855600 $Y=663340
X1323 4664 1 2 4661 DELA $T=860560 709080 1 0 $X=860560 $Y=703660
X1324 4716 1 2 4749 DELA $T=863040 668760 1 0 $X=863040 $Y=663340
X1325 5177 1 2 5154 DELA $T=937440 588120 1 0 $X=937440 $Y=582700
X1326 5095 1 2 5075 DELA $T=976500 537720 0 0 $X=976500 $Y=537340
X1327 1047 1 2 1060 DELA $T=986420 719160 0 0 $X=986420 $Y=718780
X1328 5572 1 2 5591 DELA $T=1008740 699000 0 0 $X=1008740 $Y=698620
X1329 1084 1 2 1093 DELA $T=1009980 719160 1 0 $X=1009980 $Y=713740
X1330 5540 1 2 5576 DELA $T=1011840 628440 1 0 $X=1011840 $Y=623020
X1331 4858 1 2 4881 DELA $T=1015560 709080 1 0 $X=1015560 $Y=703660
X1332 1102 1 2 1108 DELA $T=1023620 709080 1 0 $X=1023620 $Y=703660
X1333 1115 1 2 1116 DELA $T=1034160 709080 0 0 $X=1034160 $Y=708700
X1334 1138 1 2 1144 DELA $T=1068260 709080 1 0 $X=1068260 $Y=703660
X1335 1297 12 1264 2 1 4 QDFFRBN $T=231880 608280 0 180 $X=220100 $Y=602860
X1336 1300 12 1268 2 1 5 QDFFRBN $T=232500 567960 0 180 $X=220720 $Y=562540
X1337 7 11 1288 2 1 1310 QDFFRBN $T=220720 719160 1 0 $X=220720 $Y=713740
X1338 1239 12 21 2 1 14 QDFFRBN $T=221340 547800 1 0 $X=221340 $Y=542380
X1339 1306 12 1268 2 1 6 QDFFRBN $T=233120 557880 1 180 $X=221340 $Y=557500
X1340 1285 12 1268 2 1 3 QDFFRBN $T=233120 588120 0 180 $X=221340 $Y=582700
X1341 1303 12 1268 2 1 8 QDFFRBN $T=233120 598200 0 180 $X=221340 $Y=592780
X1342 1301 12 1264 2 1 9 QDFFRBN $T=233120 618360 1 180 $X=221340 $Y=617980
X1343 1250 12 1264 2 1 20 QDFFRBN $T=221340 648600 0 0 $X=221340 $Y=648220
X1344 1251 11 1288 2 1 22 QDFFRBN $T=221340 688920 0 0 $X=221340 $Y=688540
X1345 1252 11 1288 2 1 1312 QDFFRBN $T=221340 699000 1 0 $X=221340 $Y=693580
X1346 1253 11 1288 2 1 1244 QDFFRBN $T=221340 709080 1 0 $X=221340 $Y=703660
X1347 1258 12 1264 2 1 15 QDFFRBN $T=221960 638520 0 0 $X=221960 $Y=638140
X1348 1262 12 21 2 1 26 QDFFRBN $T=222580 537720 0 0 $X=222580 $Y=537340
X1349 1332 11 1288 2 1 1350 QDFFRBN $T=235600 699000 1 0 $X=235600 $Y=693580
X1350 1384 11 1288 2 1 1339 QDFFRBN $T=248620 709080 0 180 $X=236840 $Y=703660
X1351 1373 12 21 2 1 1465 QDFFRBN $T=246760 547800 1 0 $X=246760 $Y=542380
X1352 1407 11 37 2 1 1485 QDFFRBN $T=249860 709080 1 0 $X=249860 $Y=703660
X1353 1417 11 37 2 1 1409 QDFFRBN $T=250480 709080 0 0 $X=250480 $Y=708700
X1354 1461 12 1438 2 1 44 QDFFRBN $T=257300 557880 0 0 $X=257300 $Y=557500
X1355 1505 12 1438 2 1 46 QDFFRBN $T=269080 578040 1 180 $X=257300 $Y=577660
X1356 1476 12 1438 2 1 1513 QDFFRBN $T=260400 567960 1 0 $X=260400 $Y=562540
X1357 1480 12 1438 2 1 1528 QDFFRBN $T=261020 578040 1 0 $X=261020 $Y=572620
X1358 1486 12 1508 2 1 58 QDFFRBN $T=263500 628440 1 0 $X=263500 $Y=623020
X1359 1487 11 37 2 1 1545 QDFFRBN $T=263500 709080 1 0 $X=263500 $Y=703660
X1360 1546 12 1508 2 1 1491 QDFFRBN $T=276520 638520 0 180 $X=264740 $Y=633100
X1361 1503 12 1530 2 1 1564 QDFFRBN $T=266600 588120 1 0 $X=266600 $Y=582700
X1362 1506 12 1508 2 1 1576 QDFFRBN $T=267220 618360 1 0 $X=267220 $Y=612940
X1363 1517 12 1530 2 1 1580 QDFFRBN $T=269700 598200 1 0 $X=269700 $Y=592780
X1364 1519 12 1508 2 1 1531 QDFFRBN $T=270320 608280 1 0 $X=270320 $Y=602860
X1365 1542 12 1508 2 1 1578 QDFFRBN $T=274040 608280 0 0 $X=274040 $Y=607900
X1366 1598 12 1508 2 1 1509 QDFFRBN $T=288300 628440 1 180 $X=276520 $Y=628060
X1367 1563 11 1585 2 1 1547 QDFFRBN $T=277140 709080 1 0 $X=277140 $Y=703660
X1368 1569 11 37 2 1 56 QDFFRBN $T=279000 709080 0 0 $X=279000 $Y=708700
X1369 85 11 101 2 1 1681 QDFFRBN $T=287680 719160 0 0 $X=287680 $Y=718780
X1370 1625 12 1530 2 1 1641 QDFFRBN $T=290780 588120 0 0 $X=290780 $Y=587740
X1371 1689 11 1585 2 1 1635 QDFFRBN $T=303180 699000 1 180 $X=291400 $Y=698620
X1372 1636 11 84 2 1 1657 QDFFRBN $T=291400 719160 1 0 $X=291400 $Y=713740
X1373 1708 12 1530 2 1 1654 QDFFRBN $T=306900 588120 0 180 $X=295120 $Y=582700
X1374 1700 12 1623 2 1 1738 QDFFRBN $T=303800 638520 1 0 $X=303800 $Y=633100
X1375 1710 11 1755 2 1 1706 QDFFRBN $T=305660 668760 0 0 $X=305660 $Y=668380
X1376 1717 12 1623 2 1 1765 QDFFRBN $T=306900 588120 1 0 $X=306900 $Y=582700
X1377 1715 11 1775 2 1 1740 QDFFRBN $T=308140 668760 1 0 $X=308140 $Y=663340
X1378 1732 11 101 2 1 1697 QDFFRBN $T=319920 719160 1 180 $X=308140 $Y=718780
X1379 1831 136 1775 2 1 124 QDFFRBN $T=326120 658680 0 180 $X=314340 $Y=653260
X1380 1769 12 1809 2 1 125 QDFFRBN $T=315580 638520 1 0 $X=315580 $Y=633100
X1381 1777 12 1623 2 1 1799 QDFFRBN $T=316200 628440 1 0 $X=316200 $Y=623020
X1382 1778 11 1818 2 1 1810 QDFFRBN $T=316820 678840 1 0 $X=316820 $Y=673420
X1383 1779 11 1818 2 1 123 QDFFRBN $T=319300 719160 1 0 $X=319300 $Y=713740
X1384 1792 12 121 2 1 1816 QDFFRBN $T=319920 578040 1 0 $X=319920 $Y=572620
X1385 1798 11 1818 2 1 132 QDFFRBN $T=321160 699000 0 0 $X=321160 $Y=698620
X1386 1753 12 1809 2 1 1730 QDFFRBN $T=321780 578040 0 0 $X=321780 $Y=577660
X1387 1819 11 1818 2 1 1864 QDFFRBN $T=324880 668760 0 0 $X=324880 $Y=668380
X1388 1821 12 1809 2 1 1863 QDFFRBN $T=325500 588120 0 0 $X=325500 $Y=587740
X1389 1839 12 1809 2 1 141 QDFFRBN $T=329840 628440 0 0 $X=329840 $Y=628060
X1390 1888 136 1775 2 1 1844 QDFFRBN $T=342860 668760 0 180 $X=331080 $Y=663340
X1391 1848 12 1809 2 1 1840 QDFFRBN $T=331700 618360 1 0 $X=331700 $Y=612940
X1392 1803 12 148 2 1 1842 QDFFRBN $T=332320 628440 1 0 $X=332320 $Y=623020
X1393 1924 136 1809 2 1 1871 QDFFRBN $T=349680 588120 0 180 $X=337900 $Y=582700
X1394 1872 136 1775 2 1 138 QDFFRBN $T=339760 658680 1 0 $X=339760 $Y=653260
X1395 1909 136 1775 2 1 152 QDFFRBN $T=344720 648600 0 0 $X=344720 $Y=648220
X1396 1929 136 1967 2 1 1979 QDFFRBN $T=347200 668760 1 0 $X=347200 $Y=663340
X1397 1952 136 1984 2 1 1969 QDFFRBN $T=352160 588120 1 0 $X=352160 $Y=582700
X1398 1953 136 1966 2 1 1925 QDFFRBN $T=352160 618360 1 0 $X=352160 $Y=612940
X1399 1943 136 1966 2 1 159 QDFFRBN $T=352780 638520 1 0 $X=352780 $Y=633100
X1400 1921 136 1984 2 1 165 QDFFRBN $T=354020 628440 1 0 $X=354020 $Y=623020
X1401 2004 136 1967 2 1 1869 QDFFRBN $T=365800 658680 0 180 $X=354020 $Y=653260
X1402 1944 136 1961 2 1 157 QDFFRBN $T=354640 638520 0 0 $X=354640 $Y=638140
X1403 1972 136 1966 2 1 2018 QDFFRBN $T=355880 648600 1 0 $X=355880 $Y=643180
X1404 1989 136 1966 2 1 2045 QDFFRBN $T=360840 648600 0 0 $X=360840 $Y=648220
X1405 2002 136 1984 2 1 1997 QDFFRBN $T=363320 578040 0 0 $X=363320 $Y=577660
X1406 2010 136 1961 2 1 2058 QDFFRBN $T=364560 638520 1 0 $X=364560 $Y=633100
X1407 2072 136 1961 2 1 1991 QDFFRBN $T=377580 628440 0 180 $X=365800 $Y=623020
X1408 2027 136 1984 2 1 2066 QDFFRBN $T=367660 588120 1 0 $X=367660 $Y=582700
X1409 2054 136 1967 2 1 2019 QDFFRBN $T=380060 658680 0 180 $X=368280 $Y=653260
X1410 2013 136 1984 2 1 2016 QDFFRBN $T=370760 608280 1 0 $X=370760 $Y=602860
X1411 2025 136 1984 2 1 2081 QDFFRBN $T=371380 618360 1 0 $X=371380 $Y=612940
X1412 2073 136 2112 2 1 2129 QDFFRBN $T=375720 638520 0 0 $X=375720 $Y=638140
X1413 2074 136 2112 2 1 2135 QDFFRBN $T=375720 648600 0 0 $X=375720 $Y=648220
X1414 2077 136 1961 2 1 2131 QDFFRBN $T=376960 638520 1 0 $X=376960 $Y=633100
X1415 2079 136 2123 2 1 2107 QDFFRBN $T=377580 628440 1 0 $X=377580 $Y=623020
X1416 2087 136 2123 2 1 2014 QDFFRBN $T=378820 608280 0 0 $X=378820 $Y=607900
X1417 2115 136 2123 2 1 2133 QDFFRBN $T=383780 608280 1 0 $X=383780 $Y=602860
X1418 2140 136 2112 2 1 2173 QDFFRBN $T=388740 648600 1 0 $X=388740 $Y=643180
X1419 2144 136 2190 2 1 201 QDFFRBN $T=389360 588120 0 0 $X=389360 $Y=587740
X1420 2146 136 2123 2 1 2195 QDFFRBN $T=389360 628440 1 0 $X=389360 $Y=623020
X1421 2151 136 2112 2 1 2194 QDFFRBN $T=389980 638520 0 0 $X=389980 $Y=638140
X1422 2114 136 2190 2 1 196 QDFFRBN $T=392460 588120 1 0 $X=392460 $Y=582700
X1423 2170 136 2212 2 1 2179 QDFFRBN $T=393080 618360 1 0 $X=393080 $Y=612940
X1424 2185 136 2112 2 1 2186 QDFFRBN $T=395560 648600 0 0 $X=395560 $Y=648220
X1425 2110 136 2212 2 1 2172 QDFFRBN $T=396180 598200 0 0 $X=396180 $Y=597820
X1426 2191 136 2212 2 1 2216 QDFFRBN $T=402380 608280 0 0 $X=402380 $Y=607900
X1427 2229 136 2253 2 1 2243 QDFFRBN $T=403620 638520 1 0 $X=403620 $Y=633100
X1428 2136 136 2253 2 1 2219 QDFFRBN $T=404240 628440 0 0 $X=404240 $Y=628060
X1429 2251 136 2212 2 1 2236 QDFFRBN $T=407960 598200 0 0 $X=407960 $Y=597820
X1430 2223 136 2190 2 1 2312 QDFFRBN $T=408580 588120 0 0 $X=408580 $Y=587740
X1431 2309 136 2253 2 1 2252 QDFFRBN $T=420360 638520 1 180 $X=408580 $Y=638140
X1432 2308 136 2123 2 1 2257 QDFFRBN $T=421600 608280 0 180 $X=409820 $Y=602860
X1433 2267 136 2190 2 1 2357 QDFFRBN $T=411680 588120 1 0 $X=411680 $Y=582700
X1434 2193 136 2212 2 1 2271 QDFFRBN $T=412920 618360 0 0 $X=412920 $Y=617980
X1435 2315 136 2253 2 1 2305 QDFFRBN $T=418500 638520 1 0 $X=418500 $Y=633100
X1436 2304 136 2385 2 1 2350 QDFFRBN $T=421600 598200 0 0 $X=421600 $Y=597820
X1437 2328 136 2385 2 1 2351 QDFFRBN $T=422840 618360 1 0 $X=422840 $Y=612940
X1438 2341 136 2385 2 1 2389 QDFFRBN $T=423460 608280 1 0 $X=423460 $Y=602860
X1439 2347 136 2253 2 1 2334 QDFFRBN $T=424700 618360 0 0 $X=424700 $Y=617980
X1440 2360 136 2190 2 1 2388 QDFFRBN $T=425940 588120 1 0 $X=425940 $Y=582700
X1441 2376 136 2253 2 1 2370 QDFFRBN $T=427800 628440 1 0 $X=427800 $Y=623020
X1442 2399 136 2385 2 1 2356 QDFFRBN $T=432140 608280 0 0 $X=432140 $Y=607900
X1443 2423 136 259 2 1 238 QDFFRBN $T=442680 557880 1 0 $X=442680 $Y=552460
X1444 2494 136 2410 2 1 2349 QDFFRBN $T=454460 578040 0 180 $X=442680 $Y=572620
X1445 2461 136 2410 2 1 2513 QDFFRBN $T=442680 578040 0 0 $X=442680 $Y=577660
X1446 2462 136 2410 2 1 2413 QDFFRBN $T=442680 588120 0 0 $X=442680 $Y=587740
X1447 2478 136 2410 2 1 2359 QDFFRBN $T=455080 567960 0 180 $X=443300 $Y=562540
X1448 2711 311 301 2 1 292 QDFFRBN $T=489180 709080 1 180 $X=477400 $Y=708700
X1449 2756 311 301 2 1 2669 QDFFRBN $T=491660 719160 0 180 $X=479880 $Y=713740
X1450 2735 311 2788 2 1 2811 QDFFRBN $T=491040 709080 1 0 $X=491040 $Y=703660
X1451 334 311 301 2 1 320 QDFFRBN $T=503440 719160 1 180 $X=491660 $Y=718780
X1452 2757 311 2788 2 1 2818 QDFFRBN $T=493520 719160 1 0 $X=493520 $Y=713740
X1453 2796 311 2788 2 1 2795 QDFFRBN $T=500960 699000 0 0 $X=500960 $Y=698620
X1454 2819 311 2788 2 1 2886 QDFFRBN $T=505300 719160 0 0 $X=505300 $Y=718780
X1455 2936 311 2788 2 1 2874 QDFFRBN $T=527000 709080 0 180 $X=515220 $Y=703660
X1456 2988 311 2788 2 1 2934 QDFFRBN $T=536920 699000 0 180 $X=525140 $Y=693580
X1457 2950 385 393 2 1 2942 QDFFRBN $T=528240 537720 0 0 $X=528240 $Y=537340
X1458 2969 311 384 2 1 2965 QDFFRBN $T=531960 719160 1 0 $X=531960 $Y=713740
X1459 3046 311 3017 2 1 2984 QDFFRBN $T=547460 699000 1 180 $X=535680 $Y=698620
X1460 3065 311 3017 2 1 3016 QDFFRBN $T=550560 699000 0 180 $X=538780 $Y=693580
X1461 3003 385 393 2 1 2937 QDFFRBN $T=551180 557880 1 180 $X=539400 $Y=557500
X1462 398 385 393 2 1 295 QDFFRBN $T=540020 537720 0 0 $X=540020 $Y=537340
X1463 3097 311 384 2 1 412 QDFFRBN $T=559240 719160 1 180 $X=547460 $Y=718780
X1464 3126 311 3017 2 1 3093 QDFFRBN $T=565440 699000 0 180 $X=553660 $Y=693580
X1465 3140 311 3017 2 1 2681 QDFFRBN $T=566060 688920 0 180 $X=554280 $Y=683500
X1466 3128 311 459 2 1 466 QDFFRBN $T=561100 719160 0 0 $X=561100 $Y=718780
X1467 3134 311 3171 2 1 2949 QDFFRBN $T=562340 688920 0 0 $X=562340 $Y=688540
X1468 3231 311 1967 2 1 2948 QDFFRBN $T=580320 678840 0 180 $X=568540 $Y=673420
X1469 3165 311 3171 2 1 2830 QDFFRBN $T=569160 688920 1 0 $X=569160 $Y=683500
X1470 3210 311 3171 2 1 460 QDFFRBN $T=581560 709080 1 180 $X=569780 $Y=708700
X1471 492 311 459 2 1 472 QDFFRBN $T=585900 719160 1 180 $X=574120 $Y=718780
X1472 3236 311 3171 2 1 2767 QDFFRBN $T=587140 678840 1 180 $X=575360 $Y=678460
X1473 3257 311 3171 2 1 3204 QDFFRBN $T=588380 709080 0 180 $X=576600 $Y=703660
X1474 3311 3292 1967 2 1 2851 QDFFRBN $T=596440 668760 0 180 $X=584660 $Y=663340
X1475 3273 311 459 2 1 491 QDFFRBN $T=599540 719160 1 180 $X=587760 $Y=718780
X1476 3277 311 3310 2 1 2743 QDFFRBN $T=590240 678840 0 0 $X=590240 $Y=678460
X1477 3325 3292 1967 2 1 3295 QDFFRBN $T=608840 658680 0 180 $X=597060 $Y=653260
X1478 3314 3292 3353 2 1 3374 QDFFRBN $T=598920 608280 1 0 $X=598920 $Y=602860
X1479 3315 3292 3353 2 1 3303 QDFFRBN $T=598920 618360 1 0 $X=598920 $Y=612940
X1480 3317 311 3354 2 1 558 QDFFRBN $T=598920 709080 1 0 $X=598920 $Y=703660
X1481 3331 3292 3373 2 1 3040 QDFFRBN $T=602020 648600 1 0 $X=602020 $Y=643180
X1482 3333 3292 3353 2 1 3390 QDFFRBN $T=602640 598200 0 0 $X=602640 $Y=597820
X1483 3409 569 3354 2 1 3343 QDFFRBN $T=616280 678840 1 180 $X=604500 $Y=678460
X1484 3397 569 3354 2 1 542 QDFFRBN $T=616280 688920 0 180 $X=604500 $Y=683500
X1485 2901 3292 3310 2 1 3413 QDFFRBN $T=605740 668760 0 0 $X=605740 $Y=668380
X1486 3357 3292 3310 2 1 2883 QDFFRBN $T=606980 658680 0 0 $X=606980 $Y=658300
X1487 3417 569 3354 2 1 40 QDFFRBN $T=618760 688920 1 180 $X=606980 $Y=688540
X1488 3386 3292 3353 2 1 3406 QDFFRBN $T=613180 608280 1 0 $X=613180 $Y=602860
X1489 3387 569 588 2 1 2885 QDFFRBN $T=613180 709080 0 0 $X=613180 $Y=708700
X1490 3405 3292 3373 2 1 3463 QDFFRBN $T=615660 648600 0 0 $X=615660 $Y=648220
X1491 3407 569 588 2 1 554 QDFFRBN $T=615660 719160 1 0 $X=615660 $Y=713740
X1492 2945 3292 3310 2 1 3457 QDFFRBN $T=617520 658680 1 0 $X=617520 $Y=653260
X1493 3487 3292 3310 2 1 2925 QDFFRBN $T=631780 668760 1 180 $X=620000 $Y=668380
X1494 603 569 588 2 1 583 QDFFRBN $T=631780 719160 1 180 $X=620000 $Y=718780
X1495 3465 3292 3353 2 1 3266 QDFFRBN $T=627440 608280 1 0 $X=627440 $Y=602860
X1496 3472 3292 3499 2 1 3402 QDFFRBN $T=628680 638520 1 0 $X=628680 $Y=633100
X1497 3473 569 588 2 1 621 QDFFRBN $T=628680 709080 0 0 $X=628680 $Y=708700
X1498 3495 3292 3499 2 1 3565 QDFFRBN $T=631160 618360 0 0 $X=631160 $Y=617980
X1499 3501 3292 3518 2 1 3526 QDFFRBN $T=631780 658680 1 0 $X=631780 $Y=653260
X1500 3507 3292 3561 2 1 3559 QDFFRBN $T=633640 668760 0 0 $X=633640 $Y=668380
X1501 3524 569 3561 2 1 3533 QDFFRBN $T=635500 688920 1 0 $X=635500 $Y=683500
X1502 3534 569 3561 2 1 2798 QDFFRBN $T=637360 678840 0 0 $X=637360 $Y=678460
X1503 3536 3292 3575 2 1 3420 QDFFRBN $T=637980 628440 0 0 $X=637980 $Y=628060
X1504 3591 553 629 2 1 3528 QDFFRBN $T=651620 578040 0 180 $X=639840 $Y=572620
X1505 3550 3292 3575 2 1 3616 QDFFRBN $T=639840 598200 0 0 $X=639840 $Y=597820
X1506 3551 3292 3499 2 1 3589 QDFFRBN $T=639840 628440 1 0 $X=639840 $Y=623020
X1507 3556 3292 3499 2 1 3614 QDFFRBN $T=640460 608280 1 0 $X=640460 $Y=602860
X1508 630 569 3571 2 1 647 QDFFRBN $T=642940 709080 0 0 $X=642940 $Y=708700
X1509 3564 553 629 2 1 3557 QDFFRBN $T=655960 578040 1 180 $X=644180 $Y=577660
X1510 3583 3292 3626 2 1 3121 QDFFRBN $T=646040 638520 1 0 $X=646040 $Y=633100
X1511 3584 3292 3626 2 1 3631 QDFFRBN $T=646660 658680 1 0 $X=646660 $Y=653260
X1512 3636 3292 3561 2 1 3586 QDFFRBN $T=659060 668760 0 180 $X=647280 $Y=663340
X1513 653 569 3571 2 1 572 QDFFRBN $T=660300 719160 0 180 $X=648520 $Y=713740
X1514 3596 569 3561 2 1 3662 QDFFRBN $T=649140 688920 1 0 $X=649140 $Y=683500
X1515 3602 569 3645 2 1 3666 QDFFRBN $T=649760 699000 1 0 $X=649760 $Y=693580
X1516 3605 569 3645 2 1 3527 QDFFRBN $T=650380 699000 0 0 $X=650380 $Y=698620
X1517 3679 569 3571 2 1 642 QDFFRBN $T=664640 709080 0 180 $X=652860 $Y=703660
X1518 3629 553 3575 2 1 3698 QDFFRBN $T=654720 598200 1 0 $X=654720 $Y=592780
X1519 3634 553 3680 2 1 3449 QDFFRBN $T=655340 567960 0 0 $X=655340 $Y=567580
X1520 3632 553 3680 2 1 3649 QDFFRBN $T=655340 578040 1 0 $X=655340 $Y=572620
X1521 3637 553 3680 2 1 3336 QDFFRBN $T=655960 567960 1 0 $X=655960 $Y=562540
X1522 3640 553 3680 2 1 3393 QDFFRBN $T=656580 557880 0 0 $X=656580 $Y=557500
X1523 3646 553 629 2 1 3691 QDFFRBN $T=657820 547800 1 0 $X=657820 $Y=542380
X1524 3648 3292 3700 2 1 3682 QDFFRBN $T=658440 638520 1 0 $X=658440 $Y=633100
X1525 3656 3292 3700 2 1 3647 QDFFRBN $T=659060 628440 1 0 $X=659060 $Y=623020
X1526 3663 3292 3575 2 1 3703 QDFFRBN $T=660300 618360 0 0 $X=660300 $Y=617980
X1527 3667 3292 3626 2 1 3643 QDFFRBN $T=660300 668760 1 0 $X=660300 $Y=663340
X1528 3664 3292 3561 2 1 3696 QDFFRBN $T=660300 678840 1 0 $X=660300 $Y=673420
X1529 3668 3292 3659 2 1 3611 QDFFRBN $T=660920 648600 1 0 $X=660920 $Y=643180
X1530 3669 3292 3659 2 1 3041 QDFFRBN $T=660920 648600 0 0 $X=660920 $Y=648220
X1531 666 569 3571 2 1 404 QDFFRBN $T=674560 719160 0 180 $X=662780 $Y=713740
X1532 3684 569 3645 2 1 3719 QDFFRBN $T=663400 699000 1 0 $X=663400 $Y=693580
X1533 3689 569 3571 2 1 670 QDFFRBN $T=664020 709080 0 0 $X=664020 $Y=708700
X1534 3705 569 3747 2 1 3753 QDFFRBN $T=667120 678840 0 0 $X=667120 $Y=678460
X1535 3716 553 3755 2 1 3780 QDFFRBN $T=668980 557880 0 0 $X=668980 $Y=557500
X1536 3717 553 3757 2 1 3492 QDFFRBN $T=668980 578040 0 0 $X=668980 $Y=577660
X1537 3718 553 3757 2 1 3599 QDFFRBN $T=668980 588120 1 0 $X=668980 $Y=582700
X1538 3722 3292 3750 2 1 3770 QDFFRBN $T=669600 598200 0 0 $X=669600 $Y=597820
X1539 3727 553 3769 2 1 3735 QDFFRBN $T=670840 588120 0 0 $X=670840 $Y=587740
X1540 3731 553 672 2 1 3762 QDFFRBN $T=672080 547800 0 0 $X=672080 $Y=547420
X1541 3736 553 672 2 1 3598 QDFFRBN $T=673940 537720 0 0 $X=673940 $Y=537340
X1542 3743 569 3747 2 1 3777 QDFFRBN $T=673940 668760 1 0 $X=673940 $Y=663340
X1543 3740 3292 3700 2 1 3773 QDFFRBN $T=674560 628440 1 0 $X=674560 $Y=623020
X1544 3746 569 3747 2 1 3796 QDFFRBN $T=674560 678840 1 0 $X=674560 $Y=673420
X1545 3744 3292 3747 2 1 3790 QDFFRBN $T=675180 648600 0 0 $X=675180 $Y=648220
X1546 3749 569 3645 2 1 3112 QDFFRBN $T=675180 699000 0 0 $X=675180 $Y=698620
X1547 683 569 674 2 1 327 QDFFRBN $T=687580 719160 0 180 $X=675800 $Y=713740
X1548 3761 569 3645 2 1 599 QDFFRBN $T=677040 709080 1 0 $X=677040 $Y=703660
X1549 3766 569 3803 2 1 3805 QDFFRBN $T=677660 688920 1 0 $X=677660 $Y=683500
X1550 3816 553 672 2 1 673 QDFFRBN $T=690060 547800 0 180 $X=678280 $Y=542380
X1551 3767 3292 3806 2 1 3748 QDFFRBN $T=678280 628440 0 0 $X=678280 $Y=628060
X1552 3765 3292 3747 2 1 3582 QDFFRBN $T=680140 648600 1 0 $X=680140 $Y=643180
X1553 3785 3292 3822 2 1 3672 QDFFRBN $T=682000 618360 0 0 $X=682000 $Y=617980
X1554 3839 553 3755 2 1 3671 QDFFRBN $T=694400 557880 1 180 $X=682620 $Y=557500
X1555 3840 553 3757 2 1 3787 QDFFRBN $T=694400 567960 1 180 $X=682620 $Y=567580
X1556 3797 3292 3750 2 1 3821 QDFFRBN $T=684480 608280 1 0 $X=684480 $Y=602860
X1557 3800 3292 3769 2 1 3861 QDFFRBN $T=685100 598200 1 0 $X=685100 $Y=592780
X1558 3844 3292 3626 2 1 3815 QDFFRBN $T=699980 658680 1 180 $X=688200 $Y=658300
X1559 3853 569 3803 2 1 3779 QDFFRBN $T=699980 678840 1 180 $X=688200 $Y=678460
X1560 3819 569 674 2 1 686 QDFFRBN $T=688200 719160 1 0 $X=688200 $Y=713740
X1561 3829 553 3876 2 1 3881 QDFFRBN $T=691300 547800 0 0 $X=691300 $Y=547420
X1562 692 553 672 2 1 584 QDFFRBN $T=691920 547800 1 0 $X=691920 $Y=542380
X1563 3834 569 3880 2 1 3837 QDFFRBN $T=691920 709080 1 0 $X=691920 $Y=703660
X1564 3838 569 674 2 1 3809 QDFFRBN $T=691920 709080 0 0 $X=691920 $Y=708700
X1565 3841 553 3769 2 1 3482 QDFFRBN $T=692540 588120 1 0 $X=692540 $Y=582700
X1566 3842 3292 3700 2 1 3827 QDFFRBN $T=704320 628440 1 180 $X=692540 $Y=628060
X1567 3831 3292 3806 2 1 3793 QDFFRBN $T=705560 638520 0 180 $X=693780 $Y=633100
X1568 709 569 3880 2 1 696 QDFFRBN $T=708660 719160 1 180 $X=696880 $Y=718780
X1569 3878 553 3757 2 1 3904 QDFFRBN $T=699360 598200 1 0 $X=699360 $Y=592780
X1570 3879 3292 3806 2 1 3286 QDFFRBN $T=699360 628440 1 0 $X=699360 $Y=623020
X1571 3882 553 3876 2 1 3447 QDFFRBN $T=699980 557880 0 0 $X=699980 $Y=557500
X1572 3884 3292 3900 2 1 3898 QDFFRBN $T=699980 678840 1 0 $X=699980 $Y=673420
X1573 3894 569 3803 2 1 3864 QDFFRBN $T=711760 678840 1 180 $X=699980 $Y=678460
X1574 3932 553 3769 2 1 3887 QDFFRBN $T=713000 578040 0 180 $X=701220 $Y=572620
X1575 3891 3292 3912 2 1 3208 QDFFRBN $T=701840 648600 0 0 $X=701840 $Y=648220
X1576 3896 3292 3912 2 1 3625 QDFFRBN $T=703080 648600 1 0 $X=703080 $Y=643180
X1577 3942 569 3880 2 1 706 QDFFRBN $T=716100 709080 1 180 $X=704320 $Y=708700
X1578 717 553 3876 2 1 707 QDFFRBN $T=717340 537720 1 180 $X=705560 $Y=537340
X1579 3940 553 3876 2 1 3653 QDFFRBN $T=718580 547800 1 180 $X=706800 $Y=547420
X1580 3936 553 3757 2 1 3686 QDFFRBN $T=718580 588120 0 180 $X=706800 $Y=582700
X1581 3934 3292 3806 2 1 3907 QDFFRBN $T=719200 628440 1 180 $X=707420 $Y=628060
X1582 3937 3292 3914 2 1 3552 QDFFRBN $T=721060 608280 0 180 $X=709280 $Y=602860
X1583 3913 553 3955 2 1 3930 QDFFRBN $T=709900 567960 1 0 $X=709900 $Y=562540
X1584 712 569 711 2 1 514 QDFFRBN $T=710520 719160 0 0 $X=710520 $Y=718780
X1585 3923 553 3769 2 1 3956 QDFFRBN $T=711140 598200 1 0 $X=711140 $Y=592780
X1586 3926 569 3966 2 1 3963 QDFFRBN $T=711760 699000 1 0 $X=711760 $Y=693580
X1587 3929 3292 3900 2 1 3868 QDFFRBN $T=712380 668760 1 0 $X=712380 $Y=663340
X1588 3935 569 3944 2 1 3969 QDFFRBN $T=713620 678840 0 0 $X=713620 $Y=678460
X1589 3988 3292 3806 2 1 3938 QDFFRBN $T=726020 628440 0 180 $X=714240 $Y=623020
X1590 3947 553 3955 2 1 3976 QDFFRBN $T=715480 578040 1 0 $X=715480 $Y=572620
X1591 3948 3292 3986 2 1 3933 QDFFRBN $T=715480 638520 1 0 $X=715480 $Y=633100
X1592 3952 569 3966 2 1 3294 QDFFRBN $T=715480 699000 0 0 $X=715480 $Y=698620
X1593 3953 3292 3912 2 1 3993 QDFFRBN $T=716100 648600 1 0 $X=716100 $Y=643180
X1594 3922 569 3966 2 1 3018 QDFFRBN $T=716720 709080 1 0 $X=716720 $Y=703660
X1595 4015 553 3876 2 1 3945 QDFFRBN $T=730980 547800 1 180 $X=719200 $Y=547420
X1596 3961 553 3955 2 1 3924 QDFFRBN $T=720440 588120 1 0 $X=720440 $Y=582700
X1597 4023 3292 3914 2 1 3973 QDFFRBN $T=732840 598200 1 180 $X=721060 $Y=597820
X1598 3980 724 3912 2 1 4036 QDFFRBN $T=722300 658680 0 0 $X=722300 $Y=658300
X1599 3997 724 3900 2 1 3990 QDFFRBN $T=724780 678840 1 0 $X=724780 $Y=673420
X1600 4031 724 3944 2 1 4000 QDFFRBN $T=737800 699000 0 180 $X=726020 $Y=693580
X1601 4002 3292 3986 2 1 4003 QDFFRBN $T=726640 618360 0 0 $X=726640 $Y=617980
X1602 4010 553 4040 2 1 3970 QDFFRBN $T=727260 557880 0 0 $X=727260 $Y=557500
X1603 4057 724 3900 2 1 4001 QDFFRBN $T=739040 668760 0 180 $X=727260 $Y=663340
X1604 4038 724 3944 2 1 3999 QDFFRBN $T=739040 678840 1 180 $X=727260 $Y=678460
X1605 4059 742 3986 2 1 3301 QDFFRBN $T=739660 638520 0 180 $X=727880 $Y=633100
X1606 3034 724 3966 2 1 3995 QDFFRBN $T=739660 709080 1 180 $X=727880 $Y=708700
X1607 4064 553 4026 2 1 3906 QDFFRBN $T=742140 578040 0 180 $X=730360 $Y=572620
X1608 4032 553 4026 2 1 4092 QDFFRBN $T=732840 567960 1 0 $X=732840 $Y=562540
X1609 4033 3292 4070 2 1 4063 QDFFRBN $T=732840 598200 0 0 $X=732840 $Y=597820
X1610 4035 724 711 2 1 2976 QDFFRBN $T=746480 719160 1 180 $X=734700 $Y=718780
X1611 4044 742 3986 2 1 3154 QDFFRBN $T=735320 628440 1 0 $X=735320 $Y=623020
X1612 4054 553 4026 2 1 4045 QDFFRBN $T=736560 557880 1 0 $X=736560 $Y=552460
X1613 4058 553 4040 2 1 3341 QDFFRBN $T=737800 547800 0 0 $X=737800 $Y=547420
X1614 755 553 4040 2 1 768 QDFFRBN $T=739660 537720 0 0 $X=739660 $Y=537340
X1615 4125 742 4040 2 1 3515 QDFFRBN $T=752060 557880 1 180 $X=740280 $Y=557500
X1616 4117 724 3986 2 1 3378 QDFFRBN $T=752060 638520 1 180 $X=740280 $Y=638140
X1617 4071 724 4126 2 1 4119 QDFFRBN $T=742760 658680 0 0 $X=742760 $Y=658300
X1618 4089 724 740 2 1 4167 QDFFRBN $T=743380 719160 1 0 $X=743380 $Y=713740
X1619 4094 724 740 2 1 3560 QDFFRBN $T=744000 709080 1 0 $X=744000 $Y=703660
X1620 4096 742 3914 2 1 4136 QDFFRBN $T=744620 598200 0 0 $X=744620 $Y=597820
X1621 4099 742 4026 2 1 3710 QDFFRBN $T=745240 578040 1 0 $X=745240 $Y=572620
X1622 4100 742 4070 2 1 4141 QDFFRBN $T=745240 598200 1 0 $X=745240 $Y=592780
X1623 4101 742 4126 2 1 4128 QDFFRBN $T=745240 618360 1 0 $X=745240 $Y=612940
X1624 4102 724 4140 2 1 4158 QDFFRBN $T=745240 678840 1 0 $X=745240 $Y=673420
X1625 4103 724 4140 2 1 4160 QDFFRBN $T=745240 688920 0 0 $X=745240 $Y=688540
X1626 4105 742 4126 2 1 4137 QDFFRBN $T=745860 628440 0 0 $X=745860 $Y=628060
X1627 4109 742 4126 2 1 4162 QDFFRBN $T=746480 638520 1 0 $X=746480 $Y=633100
X1628 4171 742 4026 2 1 4114 QDFFRBN $T=759500 567960 0 180 $X=747720 $Y=562540
X1629 4121 724 4126 2 1 3259 QDFFRBN $T=748340 658680 1 0 $X=748340 $Y=653260
X1630 4120 742 4070 2 1 3455 QDFFRBN $T=750200 578040 0 0 $X=750200 $Y=577660
X1631 4187 742 776 2 1 4085 QDFFRBN $T=765080 537720 1 180 $X=753300 $Y=537340
X1632 4203 742 4040 2 1 4142 QDFFRBN $T=766320 547800 0 180 $X=754540 $Y=542380
X1633 4165 742 3914 2 1 4191 QDFFRBN $T=757020 608280 1 0 $X=757020 $Y=602860
X1634 4177 724 4140 2 1 4199 QDFFRBN $T=758260 699000 1 0 $X=758260 $Y=693580
X1635 4175 724 787 2 1 4226 QDFFRBN $T=758260 709080 1 0 $X=758260 $Y=703660
X1636 4178 742 4070 2 1 4213 QDFFRBN $T=758880 588120 1 0 $X=758880 $Y=582700
X1637 4230 742 4070 2 1 4179 QDFFRBN $T=771280 588120 1 180 $X=759500 $Y=587740
X1638 4185 742 4220 2 1 3496 QDFFRBN $T=760120 557880 0 0 $X=760120 $Y=557500
X1639 4174 742 4225 2 1 4193 QDFFRBN $T=760740 628440 0 0 $X=760740 $Y=628060
X1640 4195 742 4220 2 1 4214 QDFFRBN $T=761980 567960 1 0 $X=761980 $Y=562540
X1641 4237 724 4140 2 1 4130 QDFFRBN $T=774380 668760 1 180 $X=762600 $Y=668380
X1642 4201 742 4225 2 1 4086 QDFFRBN $T=763220 628440 1 0 $X=763220 $Y=623020
X1643 4229 724 4140 2 1 3451 QDFFRBN $T=775620 668760 0 180 $X=763840 $Y=663340
X1644 4204 742 4220 2 1 4257 QDFFRBN $T=764460 557880 1 0 $X=764460 $Y=552460
X1645 4205 724 4133 2 1 4227 QDFFRBN $T=764460 638520 0 0 $X=764460 $Y=638140
X1646 4207 724 787 2 1 4255 QDFFRBN $T=765080 719160 1 0 $X=765080 $Y=713740
X1647 4219 724 4252 2 1 3389 QDFFRBN $T=767560 688920 1 0 $X=767560 $Y=683500
X1648 4232 742 4070 2 1 4250 QDFFRBN $T=770660 588120 1 0 $X=770660 $Y=582700
X1649 4235 724 4252 2 1 3293 QDFFRBN $T=770660 688920 0 0 $X=770660 $Y=688540
X1650 4285 724 787 2 1 4234 QDFFRBN $T=782440 709080 0 180 $X=770660 $Y=703660
X1651 4238 742 4278 2 1 4277 QDFFRBN $T=771280 588120 0 0 $X=771280 $Y=587740
X1652 4239 742 4278 2 1 4274 QDFFRBN $T=771280 608280 1 0 $X=771280 $Y=602860
X1653 4244 742 4220 2 1 3639 QDFFRBN $T=771900 567960 0 0 $X=771900 $Y=567580
X1654 4245 724 4217 2 1 4300 QDFFRBN $T=772520 658680 1 0 $X=772520 $Y=653260
X1655 4259 742 4225 2 1 4127 QDFFRBN $T=775620 628440 0 0 $X=775620 $Y=628060
X1656 4262 742 4304 2 1 4296 QDFFRBN $T=776240 638520 1 0 $X=776240 $Y=633100
X1657 4292 724 4217 2 1 4256 QDFFRBN $T=788640 668760 0 180 $X=776860 $Y=663340
X1658 4269 742 811 2 1 4295 QDFFRBN $T=778100 557880 1 0 $X=778100 $Y=552460
X1659 4282 724 4252 2 1 4301 QDFFRBN $T=779340 688920 1 0 $X=779340 $Y=683500
X1660 4341 724 4252 2 1 4284 QDFFRBN $T=792360 699000 1 180 $X=780580 $Y=698620
X1661 4290 724 4333 2 1 3298 QDFFRBN $T=781200 719160 1 0 $X=781200 $Y=713740
X1662 4316 742 4225 2 1 4291 QDFFRBN $T=793600 618360 1 180 $X=781820 $Y=617980
X1663 4347 724 4252 2 1 3323 QDFFRBN $T=794220 688920 1 180 $X=782440 $Y=688540
X1664 4320 742 4220 2 1 4280 QDFFRBN $T=796080 567960 0 180 $X=784300 $Y=562540
X1665 4308 724 4217 2 1 4361 QDFFRBN $T=784920 658680 1 0 $X=784920 $Y=653260
X1666 4321 742 4278 2 1 4242 QDFFRBN $T=797940 608280 0 180 $X=786160 $Y=602860
X1667 4315 724 4333 2 1 4352 QDFFRBN $T=786160 719160 0 0 $X=786160 $Y=718780
X1668 4356 742 4220 2 1 4319 QDFFRBN $T=798560 547800 1 180 $X=786780 $Y=547420
X1669 4329 724 4304 2 1 4305 QDFFRBN $T=789260 638520 0 0 $X=789260 $Y=638140
X1670 4366 742 4278 2 1 4339 QDFFRBN $T=803520 618360 0 180 $X=791740 $Y=612940
X1671 4348 724 4390 2 1 3281 QDFFRBN $T=792360 709080 1 0 $X=792360 $Y=703660
X1672 4395 742 4365 2 1 4351 QDFFRBN $T=805380 588120 0 180 $X=793600 $Y=582700
X1673 4354 724 4390 2 1 4379 QDFFRBN $T=794220 688920 0 0 $X=794220 $Y=688540
X1674 4394 742 4365 2 1 4334 QDFFRBN $T=807240 578040 0 180 $X=795460 $Y=572620
X1675 4443 742 4393 2 1 4376 QDFFRBN $T=809720 547800 0 180 $X=797940 $Y=542380
X1676 4388 724 4333 2 1 3443 QDFFRBN $T=799800 719160 1 0 $X=799800 $Y=713740
X1677 4389 724 4333 2 1 3344 QDFFRBN $T=799800 719160 0 0 $X=799800 $Y=718780
X1678 4407 742 4278 2 1 4344 QDFFRBN $T=812200 608280 0 180 $X=800420 $Y=602860
X1679 4400 742 4393 2 1 826 QDFFRBN $T=801660 547800 0 0 $X=801660 $Y=547420
X1680 4419 724 4417 2 1 4382 QDFFRBN $T=814680 638520 1 180 $X=802900 $Y=638140
X1681 4427 724 4390 2 1 4383 QDFFRBN $T=815920 688920 0 180 $X=804140 $Y=683500
X1682 4415 724 4446 2 1 4367 QDFFRBN $T=804760 658680 1 0 $X=804760 $Y=653260
X1683 4461 837 4390 2 1 4375 QDFFRBN $T=817780 709080 0 180 $X=806000 $Y=703660
X1684 4457 742 4365 2 1 4337 QDFFRBN $T=818400 588120 0 180 $X=806620 $Y=582700
X1685 4416 742 4431 2 1 4355 QDFFRBN $T=818400 598200 0 180 $X=806620 $Y=592780
X1686 4424 724 4458 2 1 4373 QDFFRBN $T=807240 648600 1 0 $X=807240 $Y=643180
X1687 4463 839 4393 2 1 4425 QDFFRBN $T=819640 557880 1 180 $X=807860 $Y=557500
X1688 4418 839 4431 2 1 3484 QDFFRBN $T=819640 608280 1 180 $X=807860 $Y=607900
X1689 4408 839 4417 2 1 3327 QDFFRBN $T=820880 628440 0 180 $X=809100 $Y=623020
X1690 4412 742 4431 2 1 3522 QDFFRBN $T=821500 598200 1 180 $X=809720 $Y=597820
X1691 4428 839 4431 2 1 4381 QDFFRBN $T=822740 618360 0 180 $X=810960 $Y=612940
X1692 4405 839 4431 2 1 3380 QDFFRBN $T=822740 618360 1 180 $X=810960 $Y=617980
X1693 4444 742 847 2 1 852 QDFFRBN $T=812200 547800 1 0 $X=812200 $Y=542380
X1694 4426 839 4365 2 1 3476 QDFFRBN $T=824600 578040 0 180 $X=812820 $Y=572620
X1695 4448 724 4446 2 1 3523 QDFFRBN $T=812820 648600 0 0 $X=812820 $Y=648220
X1696 4453 724 4446 2 1 3461 QDFFRBN $T=814060 678840 1 0 $X=814060 $Y=673420
X1697 853 837 836 2 1 833 QDFFRBN $T=825840 719160 1 180 $X=814060 $Y=718780
X1698 4459 839 4499 2 1 4496 QDFFRBN $T=815300 567960 0 0 $X=815300 $Y=567580
X1699 4465 724 4446 2 1 3433 QDFFRBN $T=815920 688920 1 0 $X=815920 $Y=683500
X1700 4468 837 4481 2 1 4542 QDFFRBN $T=816540 699000 0 0 $X=816540 $Y=698620
X1701 4469 837 4464 2 1 4462 QDFFRBN $T=816540 719160 1 0 $X=816540 $Y=713740
X1702 4473 839 4458 2 1 4502 QDFFRBN $T=817780 628440 0 0 $X=817780 $Y=628060
X1703 4478 837 4446 2 1 4549 QDFFRBN $T=818400 658680 1 0 $X=818400 $Y=653260
X1704 4482 724 4458 2 1 4538 QDFFRBN $T=819020 638520 0 0 $X=819020 $Y=638140
X1705 4483 837 4446 2 1 4520 QDFFRBN $T=819020 668760 1 0 $X=819020 $Y=663340
X1706 4484 839 4499 2 1 4560 QDFFRBN $T=819640 578040 0 0 $X=819640 $Y=577660
X1707 4485 742 4304 2 1 4569 QDFFRBN $T=819640 598200 1 0 $X=819640 $Y=592780
X1708 4503 839 4393 2 1 4559 QDFFRBN $T=823360 557880 0 0 $X=823360 $Y=557500
X1709 4505 839 4304 2 1 4575 QDFFRBN $T=823360 608280 1 0 $X=823360 $Y=602860
X1710 4514 839 4304 2 1 4506 QDFFRBN $T=825220 618360 1 0 $X=825220 $Y=612940
X1711 4592 839 847 2 1 4518 QDFFRBN $T=837620 547800 0 180 $X=825840 $Y=542380
X1712 872 837 836 2 1 859 QDFFRBN $T=838860 719160 1 180 $X=827080 $Y=718780
X1713 4598 839 4499 2 1 4536 QDFFRBN $T=840100 578040 0 180 $X=828320 $Y=572620
X1714 4620 839 4458 2 1 4539 QDFFRBN $T=840100 648600 0 180 $X=828320 $Y=643180
X1715 4546 837 4481 2 1 4535 QDFFRBN $T=828940 688920 0 0 $X=828940 $Y=688540
X1716 4547 837 4464 2 1 4581 QDFFRBN $T=828940 719160 1 0 $X=828940 $Y=713740
X1717 4551 839 4595 2 1 875 QDFFRBN $T=829560 628440 1 0 $X=829560 $Y=623020
X1718 4614 839 847 2 1 865 QDFFRBN $T=841960 537720 1 180 $X=830180 $Y=537340
X1719 4558 839 4601 2 1 4512 QDFFRBN $T=830180 567960 1 0 $X=830180 $Y=562540
X1720 4563 837 4481 2 1 4491 QDFFRBN $T=830800 709080 1 0 $X=830800 $Y=703660
X1721 4605 837 4651 2 1 4656 QDFFRBN $T=838240 699000 0 0 $X=838240 $Y=698620
X1722 4608 839 4595 2 1 4621 QDFFRBN $T=838860 618360 1 0 $X=838860 $Y=612940
X1723 4684 837 4464 2 1 877 QDFFRBN $T=852500 719160 1 180 $X=840720 $Y=718780
X1724 4657 839 4601 2 1 4613 QDFFRBN $T=853120 557880 1 180 $X=841340 $Y=557500
X1725 4645 839 4499 2 1 4606 QDFFRBN $T=853740 578040 0 180 $X=841960 $Y=572620
X1726 882 839 4601 2 1 883 QDFFRBN $T=842580 537720 0 0 $X=842580 $Y=537340
X1727 4631 837 4651 2 1 4509 QDFFRBN $T=842580 688920 0 0 $X=842580 $Y=688540
X1728 4634 839 4458 2 1 4686 QDFFRBN $T=843200 648600 1 0 $X=843200 $Y=643180
X1729 4635 837 4651 2 1 4624 QDFFRBN $T=843200 678840 1 0 $X=843200 $Y=673420
X1730 4638 837 887 2 1 4664 QDFFRBN $T=843820 709080 0 0 $X=843820 $Y=708700
X1731 4643 839 4689 2 1 4697 QDFFRBN $T=845060 638520 1 0 $X=845060 $Y=633100
X1732 4653 839 4689 2 1 3547 QDFFRBN $T=846300 628440 0 0 $X=846300 $Y=628060
X1733 4655 839 4683 2 1 4678 QDFFRBN $T=847540 598200 1 0 $X=847540 $Y=592780
X1734 4662 837 887 2 1 4691 QDFFRBN $T=848160 719160 1 0 $X=848160 $Y=713740
X1735 4666 839 4499 2 1 4711 QDFFRBN $T=849400 578040 0 0 $X=849400 $Y=577660
X1736 4669 839 4683 2 1 4724 QDFFRBN $T=850020 608280 1 0 $X=850020 $Y=602860
X1737 4732 837 4458 2 1 4670 QDFFRBN $T=862420 648600 1 180 $X=850640 $Y=648220
X1738 4675 839 4601 2 1 4676 QDFFRBN $T=851260 557880 1 0 $X=851260 $Y=552460
X1739 4681 839 4705 2 1 903 QDFFRBN $T=851880 618360 1 0 $X=851880 $Y=612940
X1740 4746 839 4705 2 1 4688 QDFFRBN $T=864900 618360 1 180 $X=853120 $Y=617980
X1741 4740 837 4651 2 1 4693 QDFFRBN $T=865520 699000 1 180 $X=853740 $Y=698620
X1742 4726 839 4601 2 1 4696 QDFFRBN $T=867380 557880 1 180 $X=855600 $Y=557500
X1743 912 839 4601 2 1 896 QDFFRBN $T=868000 537720 1 180 $X=856220 $Y=537340
X1744 4753 837 4651 2 1 4709 QDFFRBN $T=868000 688920 1 180 $X=856220 $Y=688540
X1745 4741 837 4738 2 1 4716 QDFFRBN $T=868620 678840 1 180 $X=856840 $Y=678460
X1746 4770 839 4689 2 1 4728 QDFFRBN $T=870480 638520 0 180 $X=858700 $Y=633100
X1747 4775 839 907 2 1 4734 QDFFRBN $T=871720 567960 0 180 $X=859940 $Y=562540
X1748 4789 839 4705 2 1 4736 QDFFRBN $T=871720 628440 0 180 $X=859940 $Y=623020
X1749 4739 837 4738 2 1 4782 QDFFRBN $T=859940 658680 0 0 $X=859940 $Y=658300
X1750 4735 839 907 2 1 4677 QDFFRBN $T=872340 578040 0 180 $X=860560 $Y=572620
X1751 4785 839 907 2 1 4730 QDFFRBN $T=874820 547800 1 180 $X=863040 $Y=547420
X1752 4754 839 4705 2 1 4774 QDFFRBN $T=863660 608280 0 0 $X=863660 $Y=607900
X1753 4810 837 4778 2 1 908 QDFFRBN $T=876680 709080 1 180 $X=864900 $Y=708700
X1754 4765 839 4683 2 1 4829 QDFFRBN $T=865520 618360 1 0 $X=865520 $Y=612940
X1755 4766 837 4805 2 1 4762 QDFFRBN $T=865520 699000 0 0 $X=865520 $Y=698620
X1756 4769 837 4805 2 1 4755 QDFFRBN $T=866140 699000 1 0 $X=866140 $Y=693580
X1757 4823 839 4705 2 1 4764 QDFFRBN $T=878540 618360 1 180 $X=866760 $Y=617980
X1758 4781 839 4820 2 1 4806 QDFFRBN $T=868620 588120 1 0 $X=868620 $Y=582700
X1759 4784 839 4820 2 1 4808 QDFFRBN $T=869240 588120 0 0 $X=869240 $Y=587740
X1760 4841 839 907 2 1 4787 QDFFRBN $T=881640 537720 1 180 $X=869860 $Y=537340
X1761 4835 839 4689 2 1 4790 QDFFRBN $T=882880 638520 0 180 $X=871100 $Y=633100
X1762 4830 837 4738 2 1 4791 QDFFRBN $T=882880 678840 1 180 $X=871100 $Y=678460
X1763 4847 839 907 2 1 4794 QDFFRBN $T=883500 567960 0 180 $X=871720 $Y=562540
X1764 4797 837 4738 2 1 4859 QDFFRBN $T=871720 668760 1 0 $X=871720 $Y=663340
X1765 4792 837 4738 2 1 4793 QDFFRBN $T=871720 688920 0 0 $X=871720 $Y=688540
X1766 4801 837 4738 2 1 4845 QDFFRBN $T=872340 658680 0 0 $X=872340 $Y=658300
X1767 4867 839 4819 2 1 4798 QDFFRBN $T=885360 557880 1 180 $X=873580 $Y=557500
X1768 4873 839 4819 2 1 4807 QDFFRBN $T=885980 578040 0 180 $X=874200 $Y=572620
X1769 4814 4818 4683 2 1 4821 QDFFRBN $T=874820 608280 1 0 $X=874820 $Y=602860
X1770 923 837 4778 2 1 921 QDFFRBN $T=876060 719160 0 0 $X=876060 $Y=718780
X1771 4826 837 4778 2 1 4858 QDFFRBN $T=877300 719160 1 0 $X=877300 $Y=713740
X1772 4839 839 4683 2 1 4899 QDFFRBN $T=879160 618360 1 0 $X=879160 $Y=612940
X1773 4860 4818 4820 2 1 4914 QDFFRBN $T=882260 598200 0 0 $X=882260 $Y=597820
X1774 4864 839 4913 2 1 4894 QDFFRBN $T=882880 638520 1 0 $X=882880 $Y=633100
X1775 4874 837 4883 2 1 4893 QDFFRBN $T=884120 678840 0 0 $X=884120 $Y=678460
X1776 4876 839 4819 2 1 4800 QDFFRBN $T=897140 567960 0 180 $X=885360 $Y=562540
X1777 4939 837 4902 2 1 4882 QDFFRBN $T=897760 668760 0 180 $X=885980 $Y=663340
X1778 4922 837 4883 2 1 4834 QDFFRBN $T=898380 688920 1 180 $X=886600 $Y=688540
X1779 4891 839 4935 2 1 944 QDFFRBN $T=887220 537720 0 0 $X=887220 $Y=537340
X1780 4892 839 4935 2 1 4954 QDFFRBN $T=887220 557880 0 0 $X=887220 $Y=557500
X1781 4866 839 4913 2 1 4780 QDFFRBN $T=887840 648600 1 0 $X=887840 $Y=643180
X1782 4921 837 4902 2 1 4885 QDFFRBN $T=899620 658680 0 180 $X=887840 $Y=653260
X1783 4901 839 4819 2 1 948 QDFFRBN $T=888460 578040 1 0 $X=888460 $Y=572620
X1784 4911 837 4883 2 1 4842 QDFFRBN $T=890320 699000 1 0 $X=890320 $Y=693580
X1785 4918 839 4819 2 1 955 QDFFRBN $T=891560 567960 0 0 $X=891560 $Y=567580
X1786 4968 4818 4820 2 1 4920 QDFFRBN $T=903960 618360 0 180 $X=892180 $Y=612940
X1787 4924 839 4819 2 1 953 QDFFRBN $T=892800 547800 1 0 $X=892800 $Y=542380
X1788 4923 4818 4929 2 1 4862 QDFFRBN $T=893420 628440 1 0 $X=893420 $Y=623020
X1789 4931 4818 4929 2 1 4956 QDFFRBN $T=894040 598200 0 0 $X=894040 $Y=597820
X1790 4932 4818 4974 2 1 4832 QDFFRBN $T=894660 638520 1 0 $X=894660 $Y=633100
X1791 4937 837 4979 2 1 4971 QDFFRBN $T=895280 709080 1 0 $X=895280 $Y=703660
X1792 4941 837 4979 2 1 952 QDFFRBN $T=895900 719160 1 0 $X=895900 $Y=713740
X1793 4945 4818 4929 2 1 5020 QDFFRBN $T=897140 588120 0 0 $X=897140 $Y=587740
X1794 4948 837 4902 2 1 4962 QDFFRBN $T=897760 668760 0 0 $X=897760 $Y=668380
X1795 5027 4818 4929 2 1 4953 QDFFRBN $T=911400 598200 0 180 $X=899620 $Y=592780
X1796 4986 4818 5039 2 1 5058 QDFFRBN $T=904580 588120 1 0 $X=904580 $Y=582700
X1797 4999 4818 4974 2 1 5068 QDFFRBN $T=906440 618360 0 0 $X=906440 $Y=617980
X1798 5032 969 4935 2 1 5001 QDFFRBN $T=918840 547800 0 180 $X=907060 $Y=542380
X1799 4996 4818 4913 2 1 5014 QDFFRBN $T=907060 628440 1 0 $X=907060 $Y=623020
X1800 5006 4818 4913 2 1 4802 QDFFRBN $T=907060 648600 1 0 $X=907060 $Y=643180
X1801 5049 837 964 2 1 5004 QDFFRBN $T=918840 719160 1 180 $X=907060 $Y=718780
X1802 5066 969 4935 2 1 5008 QDFFRBN $T=919460 557880 0 180 $X=907680 $Y=552460
X1803 5059 837 4870 2 1 5012 QDFFRBN $T=919460 688920 1 180 $X=907680 $Y=688540
X1804 4985 837 4870 2 1 4951 QDFFRBN $T=919460 699000 0 180 $X=907680 $Y=693580
X1805 5070 4818 4974 2 1 5015 QDFFRBN $T=920080 638520 0 180 $X=908300 $Y=633100
X1806 5072 970 5035 2 1 5017 QDFFRBN $T=920700 678840 0 180 $X=908920 $Y=673420
X1807 5052 970 4979 2 1 5013 QDFFRBN $T=920700 709080 0 180 $X=908920 $Y=703660
X1808 5026 4818 5039 2 1 5046 QDFFRBN $T=909540 567960 0 0 $X=909540 $Y=567580
X1809 5048 970 4902 2 1 5018 QDFFRBN $T=923180 668760 1 180 $X=911400 $Y=668380
X1810 5045 4818 5039 2 1 5095 QDFFRBN $T=913260 588120 0 0 $X=913260 $Y=587740
X1811 5031 4818 5039 2 1 5040 QDFFRBN $T=913260 598200 1 0 $X=913260 $Y=592780
X1812 5099 969 962 2 1 967 QDFFRBN $T=925660 537720 1 180 $X=913880 $Y=537340
X1813 5053 837 4979 2 1 5110 QDFFRBN $T=914500 719160 1 0 $X=914500 $Y=713740
X1814 5077 4818 4974 2 1 971 QDFFRBN $T=930000 618360 1 180 $X=918220 $Y=617980
X1815 5126 4818 4974 2 1 5079 QDFFRBN $T=932480 638520 0 180 $X=920700 $Y=633100
X1816 5084 970 5133 2 1 5125 QDFFRBN $T=921320 668760 1 0 $X=921320 $Y=663340
X1817 5085 837 5035 2 1 5003 QDFFRBN $T=921320 688920 0 0 $X=921320 $Y=688540
X1818 5141 4818 5082 2 1 5087 QDFFRBN $T=933720 628440 0 180 $X=921940 $Y=623020
X1819 5092 970 5133 2 1 5163 QDFFRBN $T=923180 648600 0 0 $X=923180 $Y=648220
X1820 5094 4818 5039 2 1 5038 QDFFRBN $T=924420 567960 0 0 $X=924420 $Y=567580
X1821 5109 4818 5039 2 1 5107 QDFFRBN $T=925040 578040 0 0 $X=925040 $Y=577660
X1822 5111 970 5127 2 1 5098 QDFFRBN $T=925040 709080 1 0 $X=925040 $Y=703660
X1823 5114 969 989 2 1 5148 QDFFRBN $T=925660 537720 0 0 $X=925660 $Y=537340
X1824 5120 4818 5082 2 1 5177 QDFFRBN $T=926900 598200 0 0 $X=926900 $Y=597820
X1825 5169 969 5137 2 1 973 QDFFRBN $T=939300 557880 1 180 $X=927520 $Y=557500
X1826 5176 970 5133 2 1 5116 QDFFRBN $T=939300 668760 1 180 $X=927520 $Y=668380
X1827 994 970 4979 2 1 984 QDFFRBN $T=939300 719160 1 180 $X=927520 $Y=718780
X1828 5135 970 5035 2 1 5193 QDFFRBN $T=929380 699000 1 0 $X=929380 $Y=693580
X1829 5145 4818 5082 2 1 5187 QDFFRBN $T=931860 618360 0 0 $X=931860 $Y=617980
X1830 5146 4818 5133 2 1 5157 QDFFRBN $T=931860 628440 0 0 $X=931860 $Y=628060
X1831 5223 4818 5133 2 1 5168 QDFFRBN $T=946740 648600 0 180 $X=934960 $Y=643180
X1832 5204 4818 5133 2 1 5160 QDFFRBN $T=947980 648600 1 180 $X=936200 $Y=648220
X1833 5206 970 5035 2 1 5132 QDFFRBN $T=947980 668760 0 180 $X=936200 $Y=663340
X1834 5175 970 5035 2 1 5184 QDFFRBN $T=936200 688920 0 0 $X=936200 $Y=688540
X1835 5213 969 989 2 1 993 QDFFRBN $T=949840 537720 1 180 $X=938060 $Y=537340
X1836 5208 4818 5201 2 1 5174 QDFFRBN $T=949840 578040 0 180 $X=938060 $Y=572620
X1837 5248 4818 5201 2 1 5173 QDFFRBN $T=949840 578040 1 180 $X=938060 $Y=577660
X1838 5229 4818 5201 2 1 5128 QDFFRBN $T=949840 588120 1 180 $X=938060 $Y=587740
X1839 5185 970 5239 2 1 5113 QDFFRBN $T=938060 709080 1 0 $X=938060 $Y=703660
X1840 5215 969 5137 2 1 5182 QDFFRBN $T=951700 557880 1 180 $X=939920 $Y=557500
X1841 5268 969 989 2 1 5192 QDFFRBN $T=954800 547800 1 180 $X=943020 $Y=547420
X1842 5224 970 5239 2 1 5228 QDFFRBN $T=944260 709080 0 0 $X=944260 $Y=708700
X1843 1008 970 5127 2 1 997 QDFFRBN $T=956040 719160 1 180 $X=944260 $Y=718780
X1844 5242 4818 5082 2 1 5203 QDFFRBN $T=956660 618360 1 180 $X=944880 $Y=617980
X1845 5241 970 983 2 1 5238 QDFFRBN $T=959140 719160 0 180 $X=947360 $Y=713740
X1846 5250 4818 5271 2 1 5289 QDFFRBN $T=948600 628440 1 0 $X=948600 $Y=623020
X1847 5306 4818 5277 2 1 5253 QDFFRBN $T=961000 648600 0 180 $X=949220 $Y=643180
X1848 5281 970 5255 2 1 5232 QDFFRBN $T=961620 688920 1 180 $X=949840 $Y=688540
X1849 5267 969 1009 2 1 1001 QDFFRBN $T=951080 537720 0 0 $X=951080 $Y=537340
X1850 5300 970 5277 2 1 5265 QDFFRBN $T=962860 668760 1 180 $X=951080 $Y=668380
X1851 5314 969 1009 2 1 5270 QDFFRBN $T=963480 557880 0 180 $X=951700 $Y=552460
X1852 5315 4818 5288 2 1 5251 QDFFRBN $T=963480 578040 1 180 $X=951700 $Y=577660
X1853 5252 4818 5201 2 1 5178 QDFFRBN $T=964100 588120 1 180 $X=952320 $Y=587740
X1854 5257 4818 5271 2 1 5199 QDFFRBN $T=964720 598200 0 180 $X=952940 $Y=592780
X1855 5259 4818 5201 2 1 5179 QDFFRBN $T=965340 567960 1 180 $X=953560 $Y=567580
X1856 5307 969 1009 2 1 1004 QDFFRBN $T=967820 547800 1 180 $X=956040 $Y=547420
X1857 5333 4818 5271 2 1 5302 QDFFRBN $T=970300 598200 1 180 $X=958520 $Y=597820
X1858 1021 970 5127 2 1 1015 QDFFRBN $T=970300 709080 1 180 $X=958520 $Y=708700
X1859 5298 4818 5271 2 1 5328 QDFFRBN $T=959140 618360 0 0 $X=959140 $Y=617980
X1860 5301 970 5255 2 1 5233 QDFFRBN $T=970920 688920 0 180 $X=959140 $Y=683500
X1861 1023 970 5127 2 1 1016 QDFFRBN $T=971540 719160 0 180 $X=959760 $Y=713740
X1862 5326 4818 5243 2 1 5263 QDFFRBN $T=972780 638520 0 180 $X=961000 $Y=633100
X1863 5309 970 5239 2 1 5231 QDFFRBN $T=972780 699000 0 180 $X=961000 $Y=693580
X1864 5330 4818 5288 2 1 5282 QDFFRBN $T=973400 578040 0 180 $X=961620 $Y=572620
X1865 5292 970 5239 2 1 5202 QDFFRBN $T=973400 709080 0 180 $X=961620 $Y=703660
X1866 5331 4818 5243 2 1 5316 QDFFRBN $T=974020 628440 0 180 $X=962240 $Y=623020
X1867 5334 1025 1009 2 1 1003 QDFFRBN $T=975260 557880 0 180 $X=963480 $Y=552460
X1868 5340 4818 5288 2 1 5249 QDFFRBN $T=975260 578040 1 180 $X=963480 $Y=577660
X1869 5324 970 5277 2 1 5258 QDFFRBN $T=975880 658680 0 180 $X=964100 $Y=653260
X1870 5318 969 1026 2 1 1002 QDFFRBN $T=964720 537720 0 0 $X=964720 $Y=537340
X1871 5329 970 5354 2 1 5367 QDFFRBN $T=964720 658680 0 0 $X=964720 $Y=658300
X1872 5322 970 5354 2 1 5269 QDFFRBN $T=964720 668760 0 0 $X=964720 $Y=668380
X1873 5337 970 5255 2 1 5227 QDFFRBN $T=976500 678840 1 180 $X=964720 $Y=678460
X1874 5332 4818 5364 2 1 5338 QDFFRBN $T=967200 598200 1 0 $X=967200 $Y=592780
X1875 5335 4818 5277 2 1 5381 QDFFRBN $T=967820 628440 0 0 $X=967820 $Y=628060
X1876 5339 4818 5341 2 1 5387 QDFFRBN $T=969060 567960 0 0 $X=969060 $Y=567580
X1877 5382 4818 5271 2 1 5293 QDFFRBN $T=980840 608280 0 180 $X=969060 $Y=602860
X1878 5343 969 5341 2 1 1035 QDFFRBN $T=970300 547800 0 0 $X=970300 $Y=547420
X1879 5344 970 5354 2 1 5397 QDFFRBN $T=970300 678840 1 0 $X=970300 $Y=673420
X1880 5347 970 5386 2 1 1030 QDFFRBN $T=971540 719160 1 0 $X=971540 $Y=713740
X1881 5351 4818 5388 2 1 5380 QDFFRBN $T=972160 648600 1 0 $X=972160 $Y=643180
X1882 5352 970 5354 2 1 5377 QDFFRBN $T=972160 688920 1 0 $X=972160 $Y=683500
X1883 5353 970 5386 2 1 5398 QDFFRBN $T=972160 709080 0 0 $X=972160 $Y=708700
X1884 5359 970 5386 2 1 5391 QDFFRBN $T=973400 699000 0 0 $X=973400 $Y=698620
X1885 5363 4818 5364 2 1 5432 QDFFRBN $T=974640 608280 0 0 $X=974640 $Y=607900
X1886 5366 4818 5341 2 1 5404 QDFFRBN $T=975260 578040 0 0 $X=975260 $Y=577660
X1887 5373 4818 5421 2 1 5409 QDFFRBN $T=977120 648600 0 0 $X=977120 $Y=648220
X1888 5452 4818 5364 2 1 5384 QDFFRBN $T=991380 618360 0 180 $X=979600 $Y=612940
X1889 5395 1025 5341 2 1 1065 QDFFRBN $T=980220 557880 0 0 $X=980220 $Y=557500
X1890 5411 4818 5364 2 1 5476 QDFFRBN $T=983320 598200 1 0 $X=983320 $Y=592780
X1891 5399 4818 5364 2 1 5342 QDFFRBN $T=983940 608280 1 0 $X=983940 $Y=602860
X1892 5405 4818 5449 2 1 5487 QDFFRBN $T=983940 638520 0 0 $X=983940 $Y=638140
X1893 5418 970 5474 2 1 5472 QDFFRBN $T=984560 688920 1 0 $X=984560 $Y=683500
X1894 5489 4818 5449 2 1 5431 QDFFRBN $T=998200 648600 0 180 $X=986420 $Y=643180
X1895 5434 970 5386 2 1 5462 QDFFRBN $T=986420 699000 1 0 $X=986420 $Y=693580
X1896 5463 970 5386 2 1 5447 QDFFRBN $T=1000680 709080 1 180 $X=988900 $Y=708700
X1897 5528 970 5354 2 1 5468 QDFFRBN $T=1003780 678840 0 180 $X=992000 $Y=673420
X1898 5475 1025 5517 2 1 5438 QDFFRBN $T=992620 578040 1 0 $X=992620 $Y=572620
X1899 5480 4818 5449 2 1 5515 QDFFRBN $T=993860 618360 1 0 $X=993860 $Y=612940
X1900 5484 1025 5517 2 1 1080 QDFFRBN $T=995720 567960 0 0 $X=995720 $Y=567580
X1901 5493 1025 5517 2 1 5410 QDFFRBN $T=996340 567960 1 0 $X=996340 $Y=562540
X1902 5495 4818 5388 2 1 5509 QDFFRBN $T=996340 618360 0 0 $X=996340 $Y=617980
X1903 5501 970 5474 2 1 5550 QDFFRBN $T=996960 688920 1 0 $X=996960 $Y=683500
X1904 1078 970 5474 2 1 1084 QDFFRBN $T=996960 719160 0 0 $X=996960 $Y=718780
X1905 1071 1025 1059 2 1 1079 QDFFRBN $T=1009980 537720 1 180 $X=998200 $Y=537340
X1906 5507 970 5474 2 1 5533 QDFFRBN $T=998200 709080 1 0 $X=998200 $Y=703660
X1907 5508 970 5474 2 1 5562 QDFFRBN $T=998200 719160 1 0 $X=998200 $Y=713740
X1908 5510 4818 5388 2 1 5530 QDFFRBN $T=998820 638520 0 0 $X=998820 $Y=638140
X1909 5564 1025 1059 2 1 5514 QDFFRBN $T=1011840 547800 0 180 $X=1000060 $Y=542380
X1910 5556 5560 5421 2 1 5500 QDFFRBN $T=1012460 648600 0 180 $X=1000680 $Y=643180
X1911 5536 1025 5456 2 1 5558 QDFFRBN $T=1003160 578040 0 0 $X=1003160 $Y=577660
X1912 5596 4818 5388 2 1 5540 QDFFRBN $T=1015560 628440 1 180 $X=1003780 $Y=628060
X1913 5546 4818 5584 2 1 5570 QDFFRBN $T=1005020 608280 0 0 $X=1005020 $Y=607900
X1914 5551 5560 5575 2 1 5600 QDFFRBN $T=1005640 598200 1 0 $X=1005640 $Y=592780
X1915 5552 5560 5421 2 1 5548 QDFFRBN $T=1005640 658680 1 0 $X=1005640 $Y=653260
X1916 5553 970 5354 2 1 5594 QDFFRBN $T=1005640 678840 1 0 $X=1005640 $Y=673420
X1917 5624 5560 5575 2 1 5555 QDFFRBN $T=1018040 598200 1 180 $X=1006260 $Y=597820
X1918 5563 970 5616 2 1 5572 QDFFRBN $T=1007500 688920 0 0 $X=1007500 $Y=688540
X1919 5587 1025 5517 2 1 5583 QDFFRBN $T=1010600 567960 1 0 $X=1010600 $Y=562540
X1920 5593 4818 5421 2 1 5655 QDFFRBN $T=1012460 638520 0 0 $X=1012460 $Y=638140
X1921 5618 1025 1059 2 1 5588 QDFFRBN $T=1024860 547800 0 180 $X=1013080 $Y=542380
X1922 5662 1098 5611 2 1 5602 QDFFRBN $T=1025480 699000 1 180 $X=1013700 $Y=698620
X1923 5606 5560 5584 2 1 5698 QDFFRBN $T=1014320 618360 1 0 $X=1014320 $Y=612940
X1924 5613 970 5616 2 1 5634 QDFFRBN $T=1014940 688920 1 0 $X=1014940 $Y=683500
X1925 5639 5560 5584 2 1 5615 QDFFRBN $T=1027340 648600 0 180 $X=1015560 $Y=643180
X1926 5617 970 5611 2 1 5628 QDFFRBN $T=1015560 719160 1 0 $X=1015560 $Y=713740
X1927 5690 1025 5575 2 1 5599 QDFFRBN $T=1028580 578040 1 180 $X=1016800 $Y=577660
X1928 5621 1025 5671 2 1 1089 QDFFRBN $T=1017420 547800 0 0 $X=1017420 $Y=547420
X1929 5653 1025 5517 2 1 5565 QDFFRBN $T=1029200 567960 1 180 $X=1017420 $Y=567580
X1930 5676 5560 5421 2 1 5640 QDFFRBN $T=1031060 658680 0 180 $X=1019280 $Y=653260
X1931 5656 1098 5609 2 1 5641 QDFFRBN $T=1031060 678840 0 180 $X=1019280 $Y=673420
X1932 5644 5560 5575 2 1 5592 QDFFRBN $T=1031680 598200 0 180 $X=1019900 $Y=592780
X1933 5713 1098 5611 2 1 5657 QDFFRBN $T=1034160 709080 1 180 $X=1022380 $Y=708700
X1934 5661 5560 5683 2 1 5700 QDFFRBN $T=1023620 608280 0 0 $X=1023620 $Y=607900
X1935 5670 5560 5702 2 1 5689 QDFFRBN $T=1024860 598200 0 0 $X=1024860 $Y=597820
X1936 5668 5560 5584 2 1 5636 QDFFRBN $T=1024860 638520 0 0 $X=1024860 $Y=638140
X1937 5734 5560 5584 2 1 5684 QDFFRBN $T=1039740 648600 0 180 $X=1027960 $Y=643180
X1938 5740 1025 5671 2 1 5665 QDFFRBN $T=1040360 567960 0 180 $X=1028580 $Y=562540
X1939 5696 1098 5616 2 1 5678 QDFFRBN $T=1040360 688920 0 180 $X=1028580 $Y=683500
X1940 5712 1098 5616 2 1 5688 QDFFRBN $T=1040360 699000 1 180 $X=1028580 $Y=698620
X1941 5694 1025 5671 2 1 5669 QDFFRBN $T=1029200 567960 0 0 $X=1029200 $Y=567580
X1942 1114 1098 1107 2 1 1115 QDFFRBN $T=1029820 719160 0 0 $X=1029820 $Y=718780
X1943 5709 1025 5671 2 1 1105 QDFFRBN $T=1042220 557880 0 180 $X=1030440 $Y=552460
X1944 5711 1098 5609 2 1 5719 QDFFRBN $T=1031680 678840 0 0 $X=1031680 $Y=678460
X1945 5708 1098 5747 2 1 5742 QDFFRBN $T=1031680 719160 1 0 $X=1031680 $Y=713740
X1946 5722 5560 5421 2 1 5685 QDFFRBN $T=1044080 658680 0 180 $X=1032300 $Y=653260
X1947 5729 1025 1117 2 1 5679 QDFFRBN $T=1035400 537720 0 0 $X=1035400 $Y=537340
X1948 5726 5560 5765 2 1 5738 QDFFRBN $T=1035400 618360 1 0 $X=1035400 $Y=612940
X1949 5727 5560 5765 2 1 5766 QDFFRBN $T=1035400 618360 0 0 $X=1035400 $Y=617980
X1950 5787 1098 5616 2 1 5736 QDFFRBN $T=1049040 699000 0 180 $X=1037260 $Y=693580
X1951 5731 5560 5748 2 1 5454 QDFFRBN $T=1037880 638520 0 0 $X=1037880 $Y=638140
X1952 5790 1098 5748 2 1 5737 QDFFRBN $T=1049660 658680 1 180 $X=1037880 $Y=658300
X1953 5795 5560 5683 2 1 5749 QDFFRBN $T=1052760 598200 1 180 $X=1040980 $Y=597820
X1954 5809 1098 5748 2 1 5754 QDFFRBN $T=1053380 668760 1 180 $X=1041600 $Y=668380
X1955 5780 1098 5609 2 1 5753 QDFFRBN $T=1053380 688920 0 180 $X=1041600 $Y=683500
X1956 5758 1121 5702 2 1 5785 QDFFRBN $T=1042220 588120 1 0 $X=1042220 $Y=582700
X1957 5798 5560 5748 2 1 5756 QDFFRBN $T=1054000 648600 1 180 $X=1042220 $Y=648220
X1958 5803 1098 5609 2 1 5757 QDFFRBN $T=1054000 688920 1 180 $X=1042220 $Y=688540
X1959 1125 1098 5747 2 1 1119 QDFFRBN $T=1054000 719160 1 180 $X=1042220 $Y=718780
X1960 5799 5560 5683 2 1 5764 QDFFRBN $T=1055240 608280 0 180 $X=1043460 $Y=602860
X1961 5804 5560 5765 2 1 5759 QDFFRBN $T=1055860 628440 0 180 $X=1044080 $Y=623020
X1962 5820 1121 1117 2 1 5768 QDFFRBN $T=1056480 547800 0 180 $X=1044700 $Y=542380
X1963 5834 1098 5747 2 1 1122 QDFFRBN $T=1057100 719160 0 180 $X=1045320 $Y=713740
X1964 5802 5560 5765 2 1 5773 QDFFRBN $T=1049660 648600 1 0 $X=1049660 $Y=643180
X1965 5772 1121 5822 2 1 5743 QDFFRBN $T=1062060 567960 1 180 $X=1050280 $Y=567580
X1966 5808 1098 5857 2 1 5837 QDFFRBN $T=1051520 658680 0 0 $X=1051520 $Y=658300
X1967 5788 1121 5822 2 1 5814 QDFFRBN $T=1052760 567960 1 0 $X=1052760 $Y=562540
X1968 5821 5560 5863 2 1 5856 QDFFRBN $T=1052760 618360 1 0 $X=1052760 $Y=612940
X1969 5830 1121 5822 2 1 5885 QDFFRBN $T=1054000 578040 1 0 $X=1054000 $Y=572620
X1970 5831 5560 5683 2 1 5847 QDFFRBN $T=1054620 598200 0 0 $X=1054620 $Y=597820
X1971 5819 1121 5721 2 1 5843 QDFFRBN $T=1055240 588120 1 0 $X=1055240 $Y=582700
X1972 5836 1098 5865 2 1 5823 QDFFRBN $T=1055240 688920 1 0 $X=1055240 $Y=683500
X1973 5841 1098 5865 2 1 5839 QDFFRBN $T=1056480 709080 1 0 $X=1056480 $Y=703660
X1974 5902 5560 5765 2 1 5848 QDFFRBN $T=1069500 628440 0 180 $X=1057720 $Y=623020
X1975 5907 1098 5865 2 1 1132 QDFFRBN $T=1070740 719160 0 180 $X=1058960 $Y=713740
X1976 5918 1098 5865 2 1 5866 QDFFRBN $T=1073220 709080 1 180 $X=1061440 $Y=708700
X1977 5854 1098 5865 2 1 5833 QDFFRBN $T=1075080 688920 1 180 $X=1063300 $Y=688540
X1978 5917 1121 5822 2 1 5846 QDFFRBN $T=1075700 557880 0 180 $X=1063920 $Y=552460
X1979 5920 5560 5863 2 1 5879 QDFFRBN $T=1075700 648600 1 180 $X=1063920 $Y=648220
X1980 5888 1121 1143 2 1 1136 QDFFRBN $T=1064540 547800 0 0 $X=1064540 $Y=547420
X1981 5881 5560 5863 2 1 5886 QDFFRBN $T=1064540 618360 0 0 $X=1064540 $Y=617980
X1982 5882 5560 5863 2 1 5872 QDFFRBN $T=1064540 638520 1 0 $X=1064540 $Y=633100
X1983 5883 5560 5863 2 1 5939 QDFFRBN $T=1064540 648600 1 0 $X=1064540 $Y=643180
X1984 5870 1121 1143 2 1 5646 QDFFRBN $T=1065160 537720 0 0 $X=1065160 $Y=537340
X1985 5922 1121 5822 2 1 5884 QDFFRBN $T=1076940 567960 0 180 $X=1065160 $Y=562540
X1986 5889 5560 5857 2 1 5909 QDFFRBN $T=1065160 658680 0 0 $X=1065160 $Y=658300
X1987 5905 1098 5857 2 1 5929 QDFFRBN $T=1068260 688920 1 0 $X=1068260 $Y=683500
X1988 1153 1098 5936 2 1 1141 QDFFRBN $T=1083760 719160 0 180 $X=1071980 $Y=713740
X1989 5923 5560 5962 2 1 5953 QDFFRBN $T=1072600 628440 1 0 $X=1072600 $Y=623020
X1990 5924 1098 5857 2 1 5957 QDFFRBN $T=1072600 668760 0 0 $X=1072600 $Y=668380
X1991 5916 5560 5932 2 1 5927 QDFFRBN $T=1085000 588120 1 180 $X=1073220 $Y=587740
X1992 5926 5560 5932 2 1 5867 QDFFRBN $T=1085620 588120 0 180 $X=1073840 $Y=582700
X1993 5928 5560 5932 2 1 5949 QDFFRBN $T=1074460 608280 1 0 $X=1074460 $Y=602860
X1994 5984 1098 5865 2 1 5938 QDFFRBN $T=1086860 699000 0 180 $X=1075080 $Y=693580
X1995 5955 5560 5937 2 1 1147 QDFFRBN $T=1087480 578040 1 180 $X=1075700 $Y=577660
X1996 5941 5560 5975 2 1 5969 QDFFRBN $T=1075700 658680 1 0 $X=1075700 $Y=653260
X1997 5942 5560 5962 2 1 5968 QDFFRBN $T=1076320 618360 1 0 $X=1076320 $Y=612940
X1998 5944 5560 5975 2 1 5977 QDFFRBN $T=1076320 638520 0 0 $X=1076320 $Y=638140
X1999 5948 5560 5962 2 1 6000 QDFFRBN $T=1076940 638520 1 0 $X=1076940 $Y=633100
X2000 5947 1098 5989 2 1 5894 QDFFRBN $T=1077560 699000 0 0 $X=1077560 $Y=698620
X2001 5934 1121 1143 2 1 1151 QDFFRBN $T=1090580 537720 1 180 $X=1078800 $Y=537340
X2002 5954 1121 1160 2 1 5908 QDFFRBN $T=1079420 557880 0 0 $X=1079420 $Y=557500
X2003 5950 1098 5989 2 1 5978 QDFFRBN $T=1079420 709080 0 0 $X=1079420 $Y=708700
X2004 6004 1121 1143 2 1 5961 QDFFRBN $T=1092440 547800 1 180 $X=1080660 $Y=547420
X2005 5964 1121 6002 2 1 6022 QDFFRBN $T=1080660 567960 1 0 $X=1080660 $Y=562540
X2006 5967 1098 6001 2 1 5960 QDFFRBN $T=1081900 688920 1 0 $X=1081900 $Y=683500
X2007 5972 5560 5932 2 1 6009 QDFFRBN $T=1082520 608280 0 0 $X=1082520 $Y=607900
X2008 5976 5560 6002 2 1 5993 QDFFRBN $T=1083760 598200 1 0 $X=1083760 $Y=592780
X2009 5983 1098 6001 2 1 5988 QDFFRBN $T=1085000 668760 0 0 $X=1085000 $Y=668380
X2010 1158 1098 5936 2 1 1166 QDFFRBN $T=1085000 719160 1 0 $X=1085000 $Y=713740
X2011 6040 5560 1160 2 1 5986 QDFFRBN $T=1097400 578040 0 180 $X=1085620 $Y=572620
X2012 6048 1098 5857 2 1 6003 QDFFRBN $T=1100500 688920 1 180 $X=1088720 $Y=688540
X2013 6063 5560 6025 2 1 6007 QDFFRBN $T=1101740 648600 0 180 $X=1089960 $Y=643180
X2014 6018 5560 5975 2 1 5943 QDFFRBN $T=1102360 658680 0 180 $X=1090580 $Y=653260
X2015 6076 1121 1160 2 1 1163 QDFFRBN $T=1104220 537720 1 180 $X=1092440 $Y=537340
X2016 6028 1121 5937 2 1 1165 QDFFRBN $T=1093060 547800 0 0 $X=1093060 $Y=547420
X2017 6084 1098 5936 2 1 1162 QDFFRBN $T=1104840 709080 1 180 $X=1093060 $Y=708700
X2018 6036 1098 1175 2 1 6034 QDFFRBN $T=1094300 709080 1 0 $X=1094300 $Y=703660
X2019 6092 5560 6002 2 1 6021 QDFFRBN $T=1106700 598200 1 180 $X=1094920 $Y=597820
X2020 6093 5560 6002 2 1 6037 QDFFRBN $T=1107940 608280 1 180 $X=1096160 $Y=607900
X2021 6046 1098 5975 2 1 6105 QDFFRBN $T=1096160 678840 1 0 $X=1096160 $Y=673420
X2022 6047 1098 6001 2 1 6122 QDFFRBN $T=1096160 678840 0 0 $X=1096160 $Y=678460
X2023 6081 1121 1172 2 1 5990 QDFFRBN $T=1108560 567960 1 180 $X=1096780 $Y=567580
X2024 6059 5560 6025 2 1 5979 QDFFRBN $T=1109180 618360 1 180 $X=1097400 $Y=617980
X2025 6072 5560 1179 2 1 6125 QDFFRBN $T=1100500 578040 1 0 $X=1100500 $Y=572620
X2026 6087 5560 6131 2 1 6043 QDFFRBN $T=1102360 628440 1 0 $X=1102360 $Y=623020
X2027 6123 5560 6025 2 1 6073 QDFFRBN $T=1114140 638520 1 180 $X=1102360 $Y=638140
X2028 6088 5560 6131 2 1 6128 QDFFRBN $T=1102980 648600 1 0 $X=1102980 $Y=643180
X2029 6154 5560 1179 2 1 6091 QDFFRBN $T=1115380 578040 1 180 $X=1103600 $Y=577660
X2030 6095 1098 6001 2 1 6049 QDFFRBN $T=1115380 688920 1 180 $X=1103600 $Y=688540
X2031 6086 5560 6131 2 1 6139 QDFFRBN $T=1104220 648600 0 0 $X=1104220 $Y=648220
X2032 6102 1121 5937 2 1 1173 QDFFRBN $T=1119720 547800 1 180 $X=1107940 $Y=547420
X2033 6114 1121 6159 2 1 6070 QDFFRBN $T=1107940 557880 1 0 $X=1107940 $Y=552460
X2034 6130 1121 1172 2 1 6080 QDFFRBN $T=1121580 537720 1 180 $X=1109800 $Y=537340
X2035 6169 5560 6002 2 1 6107 QDFFRBN $T=1115380 598200 0 0 $X=1115380 $Y=597820
X2036 6161 5560 6181 2 1 6103 QDFFRBN $T=1116000 608280 1 0 $X=1116000 $Y=602860
X2037 6168 1098 1175 2 1 6106 QDFFRBN $T=1127780 709080 0 180 $X=1116000 $Y=703660
X2038 6183 1121 6159 2 1 6113 QDFFRBN $T=1128400 547800 0 180 $X=1116620 $Y=542380
X2039 6172 5560 6182 2 1 6142 QDFFRBN $T=1116620 578040 1 0 $X=1116620 $Y=572620
X2040 6157 5560 6182 2 1 6135 QDFFRBN $T=1116620 588120 0 0 $X=1116620 $Y=587740
X2041 6165 5560 6181 2 1 6108 QDFFRBN $T=1116620 618360 1 0 $X=1116620 $Y=612940
X2042 6177 5560 6131 2 1 6041 QDFFRBN $T=1128400 628440 0 180 $X=1116620 $Y=623020
X2043 6155 5560 6131 2 1 6082 QDFFRBN $T=1128400 638520 1 180 $X=1116620 $Y=638140
X2044 6170 5560 6131 2 1 6133 QDFFRBN $T=1128400 648600 0 180 $X=1116620 $Y=643180
X2045 6167 1098 6178 2 1 6143 QDFFRBN $T=1128400 668760 1 180 $X=1116620 $Y=668380
X2046 6175 1098 6178 2 1 6149 QDFFRBN $T=1128400 678840 1 180 $X=1116620 $Y=678460
X2047 6171 1098 6178 2 1 6071 QDFFRBN $T=1128400 688920 0 180 $X=1116620 $Y=683500
X2048 6162 1098 1175 2 1 1181 QDFFRBN $T=1128400 719160 1 180 $X=1116620 $Y=718780
X2049 6166 1121 6159 2 1 6061 QDFFRBN $T=1129020 557880 1 180 $X=1117240 $Y=557500
X2050 6152 1121 6182 2 1 1180 QDFFRBN $T=1117240 567960 1 0 $X=1117240 $Y=562540
X2051 6173 5560 6182 2 1 6160 QDFFRBN $T=1117240 578040 0 0 $X=1117240 $Y=577660
X2052 6176 5560 6181 2 1 6119 QDFFRBN $T=1117240 608280 0 0 $X=1117240 $Y=607900
X2053 6144 1098 6178 2 1 6069 QDFFRBN $T=1129020 699000 0 180 $X=1117240 $Y=693580
X2054 1992 1 2 2007 2053 2042 1233 ICV_4 $T=367660 588120 0 0 $X=367660 $Y=587740
X2055 2430 1 2 2462 2451 2494 1233 ICV_4 $T=439580 588120 1 0 $X=439580 $Y=582700
X2056 2743 1 2 2773 327 333 1233 ICV_4 $T=492280 688920 0 0 $X=492280 $Y=688540
X2057 324 1 2 332 2795 2817 1233 ICV_4 $T=496000 709080 0 0 $X=496000 $Y=708700
X2058 339 1 2 351 2818 2845 1233 ICV_4 $T=505300 709080 1 0 $X=505300 $Y=703660
X2059 2874 1 2 2917 371 2940 1233 ICV_4 $T=522040 699000 0 0 $X=522040 $Y=698620
X2060 2924 1 2 2945 2948 2970 1233 ICV_4 $T=523280 638520 0 0 $X=523280 $Y=638140
X2061 374 1 2 383 2934 2956 1233 ICV_4 $T=524520 688920 0 0 $X=524520 $Y=688540
X2062 395 1 2 401 403 410 1233 ICV_4 $T=538160 668760 0 0 $X=538160 $Y=668380
X2063 3020 1 2 3034 3040 3064 1233 ICV_4 $T=539400 628440 1 0 $X=539400 $Y=623020
X2064 429 1 2 436 438 448 1233 ICV_4 $T=557380 648600 0 0 $X=557380 $Y=648220
X2065 3112 1 2 3135 444 455 1233 ICV_4 $T=558620 678840 0 0 $X=558620 $Y=678460
X2066 501 1 2 510 514 524 1233 ICV_4 $T=589620 678840 1 0 $X=589620 $Y=673420
X2067 3298 1 2 3319 3323 3346 1233 ICV_4 $T=595820 648600 0 0 $X=595820 $Y=648220
X2068 538 1 2 3358 554 3365 1233 ICV_4 $T=603260 719160 0 0 $X=603260 $Y=718780
X2069 555 1 2 566 571 579 1233 ICV_4 $T=608840 668760 1 0 $X=608840 $Y=663340
X2070 558 1 2 3367 572 582 1233 ICV_4 $T=609460 699000 1 0 $X=609460 $Y=693580
X2071 575 1 2 585 586 594 1233 ICV_4 $T=615040 648600 1 0 $X=615040 $Y=643180
X2072 3420 1 2 3441 3443 3471 1233 ICV_4 $T=618760 618360 1 0 $X=618760 $Y=612940
X2073 3435 1 2 3456 3462 3493 1233 ICV_4 $T=621860 628440 0 0 $X=621860 $Y=628060
X2074 3482 1 2 3508 3515 3542 1233 ICV_4 $T=629920 578040 1 0 $X=629920 $Y=572620
X2075 3483 1 2 3509 614 622 1233 ICV_4 $T=629920 648600 0 0 $X=629920 $Y=648220
X2076 605 1 2 615 3526 3554 1233 ICV_4 $T=631160 678840 1 0 $X=631160 $Y=673420
X2077 3547 1 2 3566 3569 3592 1233 ICV_4 $T=639840 598200 1 0 $X=639840 $Y=592780
X2078 3559 1 2 3572 3577 3581 1233 ICV_4 $T=641080 678840 1 0 $X=641080 $Y=673420
X2079 3560 1 2 3576 3582 3606 1233 ICV_4 $T=641700 638520 0 0 $X=641700 $Y=638140
X2080 3565 1 2 3568 3589 3600 1233 ICV_4 $T=643560 618360 0 0 $X=643560 $Y=617980
X2081 3622 1 2 3628 3616 3650 1233 ICV_4 $T=654100 588120 0 0 $X=654100 $Y=587740
X2082 3639 1 2 3670 3671 3697 1233 ICV_4 $T=657200 557880 1 0 $X=657200 $Y=552460
X2083 3647 1 2 3676 3682 3677 1233 ICV_4 $T=658440 628440 0 0 $X=658440 $Y=628060
X2084 3649 1 2 3657 3686 3714 1233 ICV_4 $T=659060 578040 0 0 $X=659060 $Y=577660
X2085 654 1 2 659 647 664 1233 ICV_4 $T=661540 719160 0 0 $X=661540 $Y=718780
X2086 3735 1 2 3763 3770 3756 1233 ICV_4 $T=673940 608280 0 0 $X=673940 $Y=607900
X2087 3666 1 2 3652 670 3754 1233 ICV_4 $T=675180 699000 1 0 $X=675180 $Y=693580
X2088 3748 1 2 3751 3777 3778 1233 ICV_4 $T=675800 658680 1 0 $X=675800 $Y=653260
X2089 671 1 2 675 677 682 1233 ICV_4 $T=675800 719160 0 0 $X=675800 $Y=718780
X2090 691 1 2 697 3868 3889 1233 ICV_4 $T=692540 668760 0 0 $X=692540 $Y=668380
X2091 3861 1 2 3849 3904 3905 1233 ICV_4 $T=701840 578040 0 0 $X=701840 $Y=577660
X2092 710 1 2 714 3938 3960 1233 ICV_4 $T=709280 688920 0 0 $X=709280 $Y=688540
X2093 3887 1 2 3920 3950 3967 1233 ICV_4 $T=711140 608280 0 0 $X=711140 $Y=607900
X2094 3924 1 2 3949 3956 3959 1233 ICV_4 $T=711760 578040 0 0 $X=711760 $Y=577660
X2095 3933 1 2 3927 3886 3883 1233 ICV_4 $T=713620 648600 0 0 $X=713620 $Y=648220
X2096 3809 1 2 3804 723 726 1233 ICV_4 $T=717960 709080 0 0 $X=717960 $Y=708700
X2097 3970 1 2 3972 725 729 1233 ICV_4 $T=721060 537720 0 0 $X=721060 $Y=537340
X2098 4000 1 2 4011 3999 4018 1233 ICV_4 $T=727260 688920 1 0 $X=727260 $Y=683500
X2099 751 1 2 4084 4085 4113 1233 ICV_4 $T=738420 547800 1 0 $X=738420 $Y=542380
X2100 4119 1 2 4112 4139 4124 1233 ICV_4 $T=748340 648600 0 0 $X=748340 $Y=648220
X2101 4114 1 2 4135 4141 4143 1233 ICV_4 $T=748960 588120 1 0 $X=748960 $Y=582700
X2102 4179 1 2 4221 4242 4261 1233 ICV_4 $T=766940 618360 0 0 $X=766940 $Y=617980
X2103 4226 1 2 4197 4255 4251 1233 ICV_4 $T=770040 699000 1 0 $X=770040 $Y=693580
X2104 4250 1 2 4247 4277 4279 1233 ICV_4 $T=774380 578040 0 0 $X=774380 $Y=577660
X2105 4280 1 2 4299 4305 4330 1233 ICV_4 $T=779340 638520 0 0 $X=779340 $Y=638140
X2106 4295 1 2 4287 813 817 1233 ICV_4 $T=785540 557880 0 0 $X=785540 $Y=557500
X2107 4213 1 2 4212 4214 4236 1233 ICV_4 $T=788020 567960 0 0 $X=788020 $Y=567580
X2108 4353 1 2 4349 4319 4342 1233 ICV_4 $T=805380 628440 0 0 $X=805380 $Y=628060
X2109 4375 1 2 4432 4379 4404 1233 ICV_4 $T=807860 688920 0 0 $X=807860 $Y=688540
X2110 4496 1 2 4524 860 4529 1233 ICV_4 $T=822120 547800 0 0 $X=822120 $Y=547420
X2111 4502 1 2 4532 4538 4519 1233 ICV_4 $T=823360 638520 1 0 $X=823360 $Y=633100
X2112 4539 1 2 4607 4381 4411 1233 ICV_4 $T=843820 638520 0 0 $X=843820 $Y=638140
X2113 4676 1 2 4706 898 904 1233 ICV_4 $T=851880 547800 1 0 $X=851880 $Y=542380
X2114 4678 1 2 4682 4711 4712 1233 ICV_4 $T=851880 588120 1 0 $X=851880 $Y=582700
X2115 4619 1 2 4612 4621 4659 1233 ICV_4 $T=853120 608280 0 0 $X=853120 $Y=607900
X2116 4730 1 2 4763 915 920 1233 ICV_4 $T=863040 547800 1 0 $X=863040 $Y=542380
X2117 4802 1 2 4828 4832 4863 1233 ICV_4 $T=873580 638520 0 0 $X=873580 $Y=638140
X2118 4793 1 2 4804 929 933 1233 ICV_4 $T=877300 699000 0 0 $X=877300 $Y=698620
X2119 4862 1 2 4889 4894 4909 1233 ICV_4 $T=882880 628440 0 0 $X=882880 $Y=628060
X2120 4798 1 2 4851 943 954 1233 ICV_4 $T=892800 547800 0 0 $X=892800 $Y=547420
X2121 4807 1 2 4857 4806 4844 1233 ICV_4 $T=894040 588120 1 0 $X=894040 $Y=582700
X2122 941 1 2 951 4971 4964 1233 ICV_4 $T=897140 709080 0 0 $X=897140 $Y=708700
X2123 5003 1 2 5033 5012 5036 1233 ICV_4 $T=907060 678840 0 0 $X=907060 $Y=678460
X2124 5001 1 2 5044 5046 5047 1233 ICV_4 $T=908920 557880 0 0 $X=908920 $Y=557500
X2125 5013 1 2 5028 5004 5029 1233 ICV_4 $T=910160 709080 0 0 $X=910160 $Y=708700
X2126 5128 1 2 5152 5157 5183 1233 ICV_4 $T=928760 608280 0 0 $X=928760 $Y=607900
X2127 5160 1 2 5180 5254 5279 1233 ICV_4 $T=947980 648600 0 0 $X=947980 $Y=648220
X2128 5228 1 2 5273 5233 5287 1233 ICV_4 $T=949220 699000 1 0 $X=949220 $Y=693580
X2129 5253 1 2 5290 5014 4973 1233 ICV_4 $T=960380 638520 0 0 $X=960380 $Y=638140
X2130 5231 1 2 5291 5110 5104 1233 ICV_4 $T=960380 699000 0 0 $X=960380 $Y=698620
X2131 5134 1 2 5190 5238 5210 1233 ICV_4 $T=960380 719160 0 0 $X=960380 $Y=718780
X2132 5269 1 2 5304 5193 5189 1233 ICV_4 $T=961620 688920 0 0 $X=961620 $Y=688540
X2133 5265 1 2 5283 5227 5327 1233 ICV_4 $T=963480 668760 1 0 $X=963480 $Y=663340
X2134 5289 1 2 5276 5338 5355 1233 ICV_4 $T=964100 588120 0 0 $X=964100 $Y=587740
X2135 5328 1 2 5317 5316 5321 1233 ICV_4 $T=967200 618360 1 0 $X=967200 $Y=612940
X2136 5079 1 2 5076 5380 5401 1233 ICV_4 $T=974020 638520 0 0 $X=974020 $Y=638140
X2137 4916 1 2 4919 5249 5325 1233 ICV_4 $T=975260 557880 1 0 $X=975260 $Y=552460
X2138 1030 1 2 5349 1037 1044 1233 ICV_4 $T=976500 719160 0 0 $X=976500 $Y=718780
X2139 5404 1 2 5415 5438 5471 1233 ICV_4 $T=982700 578040 1 0 $X=982700 $Y=572620
X2140 5487 1 2 5430 5530 5531 1233 ICV_4 $T=997580 628440 1 0 $X=997580 $Y=623020
X2141 5514 1 2 5549 1083 5580 1233 ICV_4 $T=1001920 557880 1 0 $X=1001920 $Y=552460
X2142 5555 1 2 5601 5600 5567 1233 ICV_4 $T=1013700 588120 1 0 $X=1013700 $Y=582700
X2143 5548 1 2 5581 5615 5626 1233 ICV_4 $T=1019900 648600 0 0 $X=1019900 $Y=648220
X2144 5646 1 2 5666 5669 5675 1233 ICV_4 $T=1020520 557880 1 0 $X=1020520 $Y=552460
X2145 5640 1 2 5660 5685 5710 1233 ICV_4 $T=1023000 668760 1 0 $X=1023000 $Y=663340
X2146 5641 1 2 5645 5719 5723 1233 ICV_4 $T=1031680 668760 0 0 $X=1031680 $Y=668380
X2147 5684 1 2 5706 5773 5796 1233 ICV_4 $T=1039740 648600 1 0 $X=1039740 $Y=643180
X2148 5785 1 2 5783 5814 5807 1233 ICV_4 $T=1047180 578040 0 0 $X=1047180 $Y=577660
X2149 5843 1 2 5844 5867 5892 1233 ICV_4 $T=1057100 578040 0 0 $X=1057100 $Y=577660
X2150 5749 1 2 5816 5764 5779 1233 ICV_4 $T=1061440 608280 0 0 $X=1061440 $Y=607900
X2151 5839 1 2 5877 5866 5915 1233 ICV_4 $T=1061440 699000 0 0 $X=1061440 $Y=698620
X2152 5871 1 2 5903 5949 5945 1233 ICV_4 $T=1072600 598200 0 0 $X=1072600 $Y=597820
X2153 1145 1 2 1148 1149 1152 1233 ICV_4 $T=1072600 719160 0 0 $X=1072600 $Y=718780
X2154 5929 1 2 5952 5957 5956 1233 ICV_4 $T=1073840 678840 1 0 $X=1073840 $Y=673420
X2155 5943 1 2 5966 5969 5971 1233 ICV_4 $T=1077560 648600 1 0 $X=1077560 $Y=643180
X2156 5979 1 2 6006 6009 6031 1233 ICV_4 $T=1085000 598200 0 0 $X=1085000 $Y=597820
X2157 5961 1 2 5985 5885 5895 1233 ICV_4 $T=1085620 567960 0 0 $X=1085620 $Y=567580
X2158 5988 1 2 5987 5960 5997 1233 ICV_4 $T=1085620 678840 0 0 $X=1085620 $Y=678460
X2159 5993 1 2 6017 6021 6050 1233 ICV_4 $T=1087480 578040 0 0 $X=1087480 $Y=577660
X2160 6007 1 2 6026 6043 6039 1233 ICV_4 $T=1091200 638520 0 0 $X=1091200 $Y=638140
X2161 5986 1 2 6035 6061 6085 1233 ICV_4 $T=1093680 567960 1 0 $X=1093680 $Y=562540
X2162 6003 1 2 6011 1171 1176 1233 ICV_4 $T=1093680 688920 1 0 $X=1093680 $Y=683500
X2163 6073 1 2 6097 6108 6121 1233 ICV_4 $T=1105460 628440 0 0 $X=1105460 $Y=628060
X2164 6034 1 2 6083 6098 6117 1233 ICV_4 $T=1106080 709080 1 0 $X=1106080 $Y=703660
X2165 6069 1 2 6120 6122 6150 1233 ICV_4 $T=1106700 688920 1 0 $X=1106700 $Y=683500
X2166 6135 1 2 6137 5927 5893 1233 ICV_4 $T=1115380 598200 1 0 $X=1115380 $Y=592780
X2167 6107 1 2 6126 6125 6111 1233 ICV_4 $T=1115380 628440 0 0 $X=1115380 $Y=628060
X2168 5977 1 2 5992 5939 5970 1233 ICV_4 $T=1116000 648600 0 0 $X=1116000 $Y=648220
X2169 6119 1 2 6147 5968 5958 1233 ICV_4 $T=1116620 618360 0 0 $X=1116620 $Y=617980
X2170 6143 1 2 6148 6041 6158 1233 ICV_4 $T=1116620 668760 1 0 $X=1116620 $Y=663340
X2171 6160 1 2 6163 6022 6020 1233 ICV_4 $T=1118480 567960 0 0 $X=1118480 $Y=567580
X2172 6149 1 2 6156 6142 6153 1233 ICV_4 $T=1118480 678840 1 0 $X=1118480 $Y=673420
X2173 1185 1 2 1187 1162 6052 1233 ICV_4 $T=1119100 719160 1 0 $X=1119100 $Y=713740
X2174 2019 1 2 2037 2083 2074 1233 ICV_5 $T=373240 668760 1 0 $X=373240 $Y=663340
X2175 2338 1 2 2376 2284 2315 1233 ICV_5 $T=428420 628440 0 0 $X=428420 $Y=628060
X2176 291 1 2 303 2681 2708 1233 ICV_5 $T=477400 699000 0 0 $X=477400 $Y=698620
X2177 2925 1 2 2947 2949 2971 1233 ICV_5 $T=523280 658680 1 0 $X=523280 $Y=653260
X2178 431 1 2 441 443 454 1233 ICV_5 $T=558620 678840 1 0 $X=558620 $Y=673420
X2179 3154 1 2 3176 470 479 1233 ICV_5 $T=567920 618360 0 0 $X=567920 $Y=617980
X2180 3301 1 2 3322 534 546 1233 ICV_5 $T=596440 628440 0 0 $X=596440 $Y=628060
X2181 3318 1 2 3333 3341 3361 1233 ICV_5 $T=599540 557880 1 0 $X=599540 $Y=552460
X2182 529 1 2 539 543 557 1233 ICV_5 $T=599540 699000 1 0 $X=599540 $Y=693580
X2183 3370 1 2 3388 3393 3418 1233 ICV_5 $T=609460 557880 1 0 $X=609460 $Y=552460
X2184 3402 1 2 3431 3433 3453 1233 ICV_5 $T=616280 588120 1 0 $X=616280 $Y=582700
X2185 3455 1 2 3488 3492 3521 1233 ICV_5 $T=626200 588120 1 0 $X=626200 $Y=582700
X2186 3484 1 2 3517 3523 3548 1233 ICV_5 $T=630540 608280 0 0 $X=630540 $Y=607900
X2187 633 1 2 3588 3598 3620 1233 ICV_5 $T=644180 557880 0 0 $X=644180 $Y=557500
X2188 3864 1 2 3875 3753 3739 1233 ICV_5 $T=698740 688920 0 0 $X=698740 $Y=688540
X2189 4092 1 2 4087 827 828 1233 ICV_5 $T=802280 557880 1 0 $X=802280 $Y=552460
X2190 911 1 2 918 4755 4788 1233 ICV_5 $T=865520 709080 1 0 $X=865520 $Y=703660
X2191 4794 1 2 4824 4696 4694 1233 ICV_5 $T=877300 557880 1 0 $X=877300 $Y=552460
X2192 1027 1 2 1032 4728 4747 1233 ICV_5 $T=973400 709080 1 0 $X=973400 $Y=703660
X2193 6049 1 2 6116 5468 5513 1233 ICV_5 $T=1115380 688920 0 0 $X=1115380 $Y=688540
X2194 6106 1 2 6145 1186 1189 1233 ICV_5 $T=1116620 699000 0 0 $X=1116620 $Y=698620
X2195 6082 1 2 6132 6080 6109 1233 ICV_5 $T=1119100 638520 1 0 $X=1119100 $Y=633100
X2196 1467 1387 2 1 1445 1444 MUX2 $T=259780 557880 0 180 $X=255440 $Y=552460
X2197 1531 1536 2 1 1510 1491 MUX2 $T=272800 608280 1 180 $X=268460 $Y=607900
X2198 1537 1540 2 1 1565 76 MUX2 $T=274660 567960 1 0 $X=274660 $Y=562540
X2199 1589 1536 2 1 1557 1509 MUX2 $T=283340 628440 0 180 $X=279000 $Y=623020
X2200 1738 1536 2 1 1707 1580 MUX2 $T=310620 628440 0 180 $X=306280 $Y=623020
X2201 1840 1536 2 1 1825 1730 MUX2 $T=331080 618360 1 180 $X=326740 $Y=617980
X2202 160 1885 2 1 1891 1894 MUX2 $T=347200 678840 0 180 $X=342860 $Y=673420
X2203 2036 1917 2 1 2013 1905 MUX2 $T=370140 608280 0 180 $X=365800 $Y=602860
X2204 2050 2056 2 1 1972 1592 MUX2 $T=372620 648600 0 180 $X=368280 $Y=643180
X2205 2059 2056 2 1 2010 1611 MUX2 $T=373860 628440 1 180 $X=369520 $Y=628060
X2206 2055 2056 2 1 1989 1616 MUX2 $T=373240 648600 1 0 $X=373240 $Y=643180
X2207 2081 1917 2 1 1996 1863 MUX2 $T=378200 608280 1 180 $X=373860 $Y=607900
X2208 2017 2056 2 1 2072 1631 MUX2 $T=373860 628440 0 0 $X=373860 $Y=628060
X2209 2119 2056 2 1 2077 1638 MUX2 $T=385020 628440 1 180 $X=380680 $Y=628060
X2210 2129 2138 2 1 2082 125 MUX2 $T=386260 648600 0 180 $X=381920 $Y=643180
X2211 2133 1917 2 1 2104 1997 MUX2 $T=386880 598200 1 180 $X=382540 $Y=597820
X2212 2135 2138 2 1 2083 124 MUX2 $T=388740 658680 1 180 $X=384400 $Y=658300
X2213 2145 2148 2 1 2079 1720 MUX2 $T=389980 618360 0 180 $X=385640 $Y=612940
X2214 2172 1917 2 1 2091 2066 MUX2 $T=393700 598200 1 180 $X=389360 $Y=597820
X2215 2173 2138 2 1 2126 152 MUX2 $T=393700 648600 1 180 $X=389360 $Y=648220
X2216 2156 2148 2 1 2170 1604 MUX2 $T=391220 608280 0 0 $X=391220 $Y=607900
X2217 2186 2138 2 1 2158 138 MUX2 $T=396180 658680 0 180 $X=391840 $Y=653260
X2218 2233 2148 2 1 2146 2039 MUX2 $T=405480 628440 0 180 $X=401140 $Y=623020
X2219 2236 2208 2 1 2215 1969 MUX2 $T=406100 598200 0 180 $X=401760 $Y=592780
X2220 2243 2138 2 1 2202 141 MUX2 $T=406100 638520 1 180 $X=401760 $Y=638140
X2221 2271 2148 2 1 2171 58 MUX2 $T=412920 618360 1 180 $X=408580 $Y=617980
X2222 2252 2138 2 1 2272 157 MUX2 $T=416640 648600 0 180 $X=412300 $Y=643180
X2223 2283 2208 2 1 2308 1950 MUX2 $T=414160 608280 0 0 $X=414160 $Y=607900
X2224 2350 2208 2 1 2282 15 MUX2 $T=425940 588120 1 180 $X=421600 $Y=587740
X2225 2370 2298 2 1 2338 1925 MUX2 $T=427800 628440 0 180 $X=423460 $Y=623020
X2226 2356 2298 2 1 2390 201 MUX2 $T=425940 608280 0 0 $X=425940 $Y=607900
X2227 2388 2380 2 1 2358 2357 MUX2 $T=430900 578040 1 180 $X=426560 $Y=577660
X2228 2389 2208 2 1 2363 196 MUX2 $T=430900 588120 1 180 $X=426560 $Y=587740
X2229 2406 246 2 1 2451 2349 MUX2 $T=435240 578040 1 0 $X=435240 $Y=572620
X2230 2413 2380 2 1 2430 2239 MUX2 $T=435860 588120 0 0 $X=435860 $Y=587740
X2231 2440 246 2 1 2423 2424 MUX2 $T=441440 557880 1 180 $X=437100 $Y=557500
X2232 2416 246 2 1 2478 2459 MUX2 $T=438960 567960 0 0 $X=438960 $Y=567580
X2233 2496 246 2 1 258 2479 MUX2 $T=450120 547800 0 180 $X=445780 $Y=542380
X2234 2845 2839 2 1 2757 343 MUX2 $T=510880 719160 0 180 $X=506540 $Y=713740
X2235 2915 2875 2 1 2819 361 MUX2 $T=519560 719160 0 180 $X=515220 $Y=713740
X2236 2917 2875 2 1 2936 340 MUX2 $T=522040 709080 0 0 $X=522040 $Y=708700
X2237 2940 2839 2 1 372 361 MUX2 $T=527000 719160 0 180 $X=522660 $Y=713740
X2238 2956 2839 2 1 2988 390 MUX2 $T=529480 709080 1 0 $X=529480 $Y=703660
X2239 2972 389 2 1 2950 2958 MUX2 $T=534440 547800 0 180 $X=530100 $Y=542380
X2240 2964 389 2 1 3003 3012 MUX2 $T=533820 557880 0 0 $X=533820 $Y=557500
X2241 2989 389 2 1 3013 3014 MUX2 $T=535060 547800 0 0 $X=535060 $Y=547420
X2242 3029 2839 2 1 3046 408 MUX2 $T=542500 709080 0 0 $X=542500 $Y=708700
X2243 3075 2875 2 1 405 407 MUX2 $T=549940 719160 0 180 $X=545600 $Y=713740
X2244 3087 3082 2 1 3065 408 MUX2 $T=553040 709080 1 180 $X=548700 $Y=708700
X2245 3086 3082 2 1 3105 427 MUX2 $T=552420 709080 1 0 $X=552420 $Y=703660
X2246 434 432 2 1 3097 407 MUX2 $T=559240 719160 0 180 $X=554900 $Y=713740
X2247 3109 2839 2 1 3126 427 MUX2 $T=557380 709080 1 0 $X=557380 $Y=703660
X2248 3367 550 2 1 3317 548 MUX2 $T=610080 709080 1 180 $X=605740 $Y=708700
X2249 3365 3368 2 1 3407 548 MUX2 $T=608840 719160 1 0 $X=608840 $Y=713740
X2250 3554 3553 2 1 3501 608 MUX2 $T=640460 668760 0 180 $X=636120 $Y=663340
X2251 3337 602 2 1 618 620 MUX2 $T=641700 719160 1 180 $X=637360 $Y=718780
X2252 3568 3567 2 1 3495 617 MUX2 $T=644180 618360 0 180 $X=639840 $Y=612940
X2253 3581 3585 2 1 3512 608 MUX2 $T=645420 668760 0 180 $X=641080 $Y=663340
X2254 3431 3553 2 1 3472 3544 MUX2 $T=646040 648600 0 180 $X=641700 $Y=643180
X2255 3600 3595 2 1 3551 617 MUX2 $T=649140 618360 0 180 $X=644800 $Y=612940
X2256 3593 3585 2 1 3486 3544 MUX2 $T=649140 648600 1 180 $X=644800 $Y=648220
X2257 3572 3585 2 1 3507 3458 MUX2 $T=651620 668760 1 180 $X=647280 $Y=668380
X2258 3628 3567 2 1 3555 3603 MUX2 $T=654720 588120 0 180 $X=650380 $Y=582700
X2259 3441 3630 2 1 3536 3544 MUX2 $T=654720 628440 1 180 $X=650380 $Y=628060
X2260 3146 3553 2 1 3583 3627 MUX2 $T=652240 648600 1 0 $X=652240 $Y=643180
X2261 3612 3553 2 1 3636 3458 MUX2 $T=652240 668760 0 0 $X=652240 $Y=668380
X2262 3642 3595 2 1 3556 646 MUX2 $T=658440 608280 0 180 $X=654100 $Y=602860
X2263 3290 3567 2 1 3465 3624 MUX2 $T=658440 618360 0 180 $X=654100 $Y=612940
X2264 3661 3585 2 1 3584 3627 MUX2 $T=658440 648600 1 180 $X=654100 $Y=648220
X2265 3657 3595 2 1 3632 3603 MUX2 $T=659680 588120 0 180 $X=655340 $Y=582700
X2266 3650 3567 2 1 3550 646 MUX2 $T=659680 598200 1 180 $X=655340 $Y=597820
X2267 3641 3587 2 1 3679 655 MUX2 $T=657820 709080 0 0 $X=657820 $Y=708700
X2268 3690 657 2 1 3646 646 MUX2 $T=665260 537720 1 180 $X=660920 $Y=537340
X2269 3699 3695 2 1 3663 3603 MUX2 $T=667120 608280 1 180 $X=662780 $Y=607900
X2270 3592 3595 2 1 3574 3624 MUX2 $T=664640 608280 1 0 $X=664640 $Y=602860
X2271 3676 3693 2 1 3656 3603 MUX2 $T=672700 628440 1 180 $X=668360 $Y=628060
X2272 3754 3587 2 1 3689 663 MUX2 $T=675800 709080 0 180 $X=671460 $Y=703660
X2273 3781 3752 2 1 3740 3603 MUX2 $T=679520 618360 1 180 $X=675180 $Y=617980
X2274 3804 3587 2 1 3838 676 MUX2 $T=685720 709080 0 0 $X=685720 $Y=708700
X2275 3814 3630 2 1 3831 3832 MUX2 $T=688200 638520 0 0 $X=688200 $Y=638140
X2276 3823 3693 2 1 3842 3832 MUX2 $T=689440 638520 1 0 $X=689440 $Y=633100
X2277 3846 3752 2 1 3797 3624 MUX2 $T=694400 598200 1 180 $X=690060 $Y=597820
X2278 3799 3732 2 1 3853 3458 MUX2 $T=690680 688920 1 0 $X=690680 $Y=683500
X2279 695 694 2 1 3819 676 MUX2 $T=695640 719160 1 180 $X=691300 $Y=718780
X2280 3863 3824 2 1 3844 3832 MUX2 $T=697500 668760 0 180 $X=693160 $Y=663340
X2281 3866 3713 2 1 3834 3701 MUX2 $T=697500 699000 1 180 $X=693160 $Y=698620
X2282 3883 3843 2 1 3851 3832 MUX2 $T=698740 648600 1 180 $X=694400 $Y=648220
X2283 3508 3847 2 1 3841 693 MUX2 $T=701220 578040 0 180 $X=696880 $Y=572620
X2284 3872 3695 2 1 3893 3624 MUX2 $T=698740 608280 1 0 $X=698740 $Y=602860
X2285 3905 3792 2 1 3878 3888 MUX2 $T=706800 588120 1 180 $X=702460 $Y=587740
X2286 3309 3732 2 1 3952 3701 MUX2 $T=708660 699000 0 0 $X=708660 $Y=698620
X2287 3714 3776 2 1 3936 3888 MUX2 $T=710520 588120 0 0 $X=710520 $Y=587740
X2288 3889 3824 2 1 3929 3958 MUX2 $T=711140 668760 0 0 $X=711140 $Y=668380
X2289 713 3587 2 1 3942 716 MUX2 $T=711140 719160 1 0 $X=711140 $Y=713740
X2290 3927 3890 2 1 3948 3958 MUX2 $T=712380 638520 0 0 $X=712380 $Y=638140
X2291 3962 3644 2 1 3935 3562 MUX2 $T=719820 678840 0 180 $X=715480 $Y=673420
X2292 3967 3885 2 1 3928 3951 MUX2 $T=720440 618360 0 180 $X=716100 $Y=612940
X2293 3943 3843 2 1 3971 3958 MUX2 $T=716100 658680 0 0 $X=716100 $Y=658300
X2294 3965 3678 2 1 3926 3562 MUX2 $T=720440 688920 0 180 $X=716100 $Y=683500
X2295 3989 3811 2 1 3953 3951 MUX2 $T=724160 638520 1 180 $X=719820 $Y=638140
X2296 3972 3856 2 1 4010 721 MUX2 $T=721060 557880 0 0 $X=721060 $Y=557500
X2297 3960 3862 2 1 3988 3951 MUX2 $T=728500 628440 1 180 $X=724160 $Y=628060
X2298 3964 3916 2 1 4015 721 MUX2 $T=725400 557880 1 0 $X=725400 $Y=552460
X2299 3957 3916 2 1 3913 715 MUX2 $T=725400 567960 1 0 $X=725400 $Y=562540
X2300 4016 3946 2 1 4023 3951 MUX2 $T=729120 608280 1 0 $X=729120 $Y=602860
X2301 4028 3968 2 1 4002 3951 MUX2 $T=733460 618360 0 180 $X=729120 $Y=612940
X2302 4011 3918 2 1 4031 3562 MUX2 $T=729120 699000 0 0 $X=729120 $Y=698620
X2303 4014 4037 2 1 3997 655 MUX2 $T=734700 668760 1 180 $X=730360 $Y=668380
X2304 4018 3897 2 1 4038 3562 MUX2 $T=730360 688920 0 0 $X=730360 $Y=688540
X2305 3588 737 2 1 4012 715 MUX2 $T=735320 537720 1 180 $X=730980 $Y=537340
X2306 3322 4048 2 1 4059 4068 MUX2 $T=735320 648600 1 0 $X=735320 $Y=643180
X2307 3925 4042 2 1 4064 748 MUX2 $T=735940 578040 0 0 $X=735940 $Y=577660
X2308 4065 4037 2 1 3980 716 MUX2 $T=740280 658680 1 180 $X=735940 $Y=658300
X2309 4074 4075 2 1 4033 748 MUX2 $T=742140 588120 1 180 $X=737800 $Y=587740
X2310 4112 4037 2 1 4071 3284 MUX2 $T=745240 658680 0 180 $X=740900 $Y=653260
X2311 3488 4042 2 1 4120 767 MUX2 $T=742140 588120 0 0 $X=742140 $Y=587740
X2312 3176 4079 2 1 4044 4116 MUX2 $T=742760 618360 0 0 $X=742760 $Y=617980
X2313 4087 4075 2 1 4032 4115 MUX2 $T=744000 567960 0 0 $X=744000 $Y=567580
X2314 3399 4037 2 1 4117 4111 MUX2 $T=744000 648600 0 0 $X=744000 $Y=648220
X2315 4131 4095 2 1 4101 4116 MUX2 $T=752060 608280 1 180 $X=747720 $Y=607900
X2316 3542 4042 2 1 4125 4115 MUX2 $T=748340 567960 0 0 $X=748340 $Y=567580
X2317 4132 4041 2 1 4105 4116 MUX2 $T=752680 628440 0 180 $X=748340 $Y=623020
X2318 3576 4090 2 1 4094 4107 MUX2 $T=752680 699000 1 180 $X=748340 $Y=698620
X2319 4073 4042 2 1 4054 4144 MUX2 $T=749580 557880 1 0 $X=749580 $Y=552460
X2320 4138 4048 2 1 4109 4116 MUX2 $T=753920 648600 0 180 $X=749580 $Y=643180
X2321 4155 4108 2 1 4103 4107 MUX2 $T=754540 688920 0 180 $X=750200 $Y=683500
X2322 3361 4075 2 1 4058 4144 MUX2 $T=761360 557880 0 180 $X=757020 $Y=552460
X2323 4113 4042 2 1 4187 4188 MUX2 $T=757640 547800 0 0 $X=757640 $Y=547420
X2324 4192 4104 2 1 4174 4173 MUX2 $T=762600 638520 0 180 $X=758260 $Y=633100
X2325 4197 4066 2 1 4175 4107 MUX2 $T=762600 699000 1 180 $X=758260 $Y=698620
X2326 3733 4042 2 1 4099 785 MUX2 $T=758880 578040 1 0 $X=758880 $Y=572620
X2327 4118 4041 2 1 4201 4173 MUX2 $T=758880 618360 0 0 $X=758880 $Y=617980
X2328 4198 4076 2 1 4177 4107 MUX2 $T=763840 688920 0 180 $X=759500 $Y=683500
X2329 4196 4075 2 1 4203 4188 MUX2 $T=762600 547800 0 0 $X=762600 $Y=547420
X2330 3282 4048 2 1 4121 4210 MUX2 $T=762600 658680 1 0 $X=762600 $Y=653260
X2331 4212 4043 2 1 4178 785 MUX2 $T=767560 578040 0 180 $X=763220 $Y=572620
X2332 4123 4079 2 1 4200 4173 MUX2 $T=768180 608280 1 180 $X=763840 $Y=607900
X2333 4236 4095 2 1 4195 785 MUX2 $T=771900 567960 1 180 $X=767560 $Y=567580
X2334 3509 4048 2 1 4243 3284 MUX2 $T=767560 658680 1 0 $X=767560 $Y=653260
X2335 4159 4037 2 1 4237 4210 MUX2 $T=767560 678840 1 0 $X=767560 $Y=673420
X2336 4084 747 2 1 795 4188 MUX2 $T=768180 537720 0 0 $X=768180 $Y=537340
X2337 4246 4043 2 1 4204 4188 MUX2 $T=772520 547800 1 180 $X=768180 $Y=547420
X2338 4221 4043 2 1 4230 4183 MUX2 $T=768180 598200 1 0 $X=768180 $Y=592780
X2339 3478 4108 2 1 4229 4111 MUX2 $T=773760 658680 1 180 $X=769420 $Y=658300
X2340 4247 4043 2 1 4232 4115 MUX2 $T=774380 578040 1 180 $X=770040 $Y=577660
X2341 4251 4066 2 1 4207 678 MUX2 $T=775000 709080 1 180 $X=770660 $Y=708700
X2342 3670 4095 2 1 4244 4115 MUX2 $T=776860 578040 0 180 $X=772520 $Y=572620
X2343 3529 4043 2 1 4185 4144 MUX2 $T=773140 557880 0 0 $X=773140 $Y=557500
X2344 4249 4095 2 1 4275 802 MUX2 $T=774380 547800 0 0 $X=774380 $Y=547420
X2345 4279 4020 2 1 4238 4183 MUX2 $T=779340 598200 1 180 $X=775000 $Y=597820
X2346 4150 4041 2 1 4259 4265 MUX2 $T=781200 618360 1 180 $X=776860 $Y=617980
X2347 4266 4090 2 1 4285 678 MUX2 $T=776860 719160 1 0 $X=776860 $Y=713740
X2348 4268 800 2 1 809 4188 MUX2 $T=777480 537720 0 0 $X=777480 $Y=537340
X2349 4287 4095 2 1 4269 4144 MUX2 $T=781820 557880 1 180 $X=777480 $Y=557500
X2350 4271 4076 2 1 4292 678 MUX2 $T=778100 668760 0 0 $X=778100 $Y=668380
X2351 4310 4076 2 1 4282 4210 MUX2 $T=786160 678840 0 180 $X=781820 $Y=673420
X2352 3319 4066 2 1 4290 807 MUX2 $T=786780 709080 0 180 $X=782440 $Y=703660
X2353 4299 4240 2 1 4320 812 MUX2 $T=783680 567960 0 0 $X=783680 $Y=567580
X2354 4261 4240 2 1 4321 4253 MUX2 $T=783680 608280 0 0 $X=783680 $Y=607900
X2355 4289 4240 2 1 4331 4183 MUX2 $T=785540 598200 0 0 $X=785540 $Y=597820
X2356 4335 4153 2 1 4245 4253 MUX2 $T=790500 648600 1 180 $X=786160 $Y=648220
X2357 4338 4079 2 1 4316 4313 MUX2 $T=791120 618360 0 180 $X=786780 $Y=612940
X2358 4318 4090 2 1 4341 807 MUX2 $T=786780 709080 1 0 $X=786780 $Y=703660
X2359 4349 4104 2 1 4328 4325 MUX2 $T=792980 628440 1 180 $X=788640 $Y=628060
X2360 4342 4240 2 1 4356 802 MUX2 $T=791120 557880 1 0 $X=791120 $Y=552460
X2361 3346 4076 2 1 4347 796 MUX2 $T=792360 688920 1 0 $X=792360 $Y=683500
X2362 3299 4090 2 1 4348 796 MUX2 $T=792980 719160 1 0 $X=792980 $Y=713740
X2363 3493 4104 2 1 4384 4357 MUX2 $T=794220 638520 1 0 $X=794220 $Y=633100
X2364 3388 4108 2 1 4340 3284 MUX2 $T=798560 668760 1 180 $X=794220 $Y=668380
X2365 820 747 2 1 4400 812 MUX2 $T=797940 537720 0 0 $X=797940 $Y=537340
X2366 4377 4240 2 1 4394 4357 MUX2 $T=797940 567960 0 0 $X=797940 $Y=567580
X2367 4370 4240 2 1 4395 4396 MUX2 $T=797940 588120 0 0 $X=797940 $Y=587740
X2368 4386 4153 2 1 4415 4210 MUX2 $T=799800 658680 1 0 $X=799800 $Y=653260
X2369 4404 4076 2 1 4354 819 MUX2 $T=804140 688920 0 180 $X=799800 $Y=683500
X2370 3408 4041 2 1 4405 4343 MUX2 $T=800420 618360 0 0 $X=800420 $Y=617980
X2371 4380 4041 2 1 4407 4396 MUX2 $T=801040 598200 0 0 $X=801040 $Y=597820
X2372 3349 4104 2 1 4408 4068 MUX2 $T=801040 628440 0 0 $X=801040 $Y=628060
X2373 3456 4108 2 1 4413 4068 MUX2 $T=801040 678840 1 0 $X=801040 $Y=673420
X2374 4397 4153 2 1 4419 4357 MUX2 $T=801660 648600 1 0 $X=801660 $Y=643180
X2375 4401 4020 2 1 4416 4396 MUX2 $T=802280 588120 0 0 $X=802280 $Y=587740
X2376 4409 4104 2 1 4424 4210 MUX2 $T=804760 648600 0 0 $X=804760 $Y=648220
X2377 4410 4076 2 1 4427 4423 MUX2 $T=804760 678840 0 0 $X=804760 $Y=678460
X2378 3549 4079 2 1 4412 4396 MUX2 $T=809720 598200 1 180 $X=805380 $Y=597820
X2379 4411 4079 2 1 4428 4343 MUX2 $T=805380 618360 1 0 $X=805380 $Y=612940
X2380 4414 4066 2 1 4429 4423 MUX2 $T=805380 699000 0 0 $X=805380 $Y=698620
X2381 4422 4020 2 1 4436 4343 MUX2 $T=807240 567960 0 0 $X=807240 $Y=567580
X2382 3471 4090 2 1 4388 4423 MUX2 $T=811580 709080 1 180 $X=807240 $Y=708700
X2383 3506 4020 2 1 4426 812 MUX2 $T=812820 578040 0 180 $X=808480 $Y=572620
X2384 4432 4090 2 1 4461 819 MUX2 $T=810340 699000 0 0 $X=810340 $Y=698620
X2385 4435 800 2 1 4443 834 MUX2 $T=810960 537720 0 0 $X=810960 $Y=537340
X2386 4439 4020 2 1 4457 818 MUX2 $T=811580 578040 0 0 $X=811580 $Y=577660
X2387 4488 4487 2 1 4463 822 MUX2 $T=820260 557880 0 180 $X=815920 $Y=552460
X2388 854 4487 2 1 4444 834 MUX2 $T=825220 557880 0 180 $X=820880 $Y=552460
X2389 4529 4530 2 1 848 834 MUX2 $T=827700 537720 1 180 $X=823360 $Y=537340
X2390 4524 4530 2 1 4459 4343 MUX2 $T=828940 567960 0 180 $X=824600 $Y=562540
X2391 4553 4530 2 1 4503 822 MUX2 $T=830800 557880 0 180 $X=826460 $Y=552460
X2392 4565 4530 2 1 4505 4537 MUX2 $T=832660 598200 1 180 $X=828320 $Y=597820
X2393 4548 4487 2 1 4558 868 MUX2 $T=829560 567960 0 0 $X=829560 $Y=567580
X2394 4541 4487 2 1 4514 4537 MUX2 $T=833900 608280 1 180 $X=829560 $Y=607900
X2395 4532 4550 2 1 4473 4582 MUX2 $T=830800 628440 0 0 $X=830800 $Y=628060
X2396 4576 4550 2 1 4478 4557 MUX2 $T=835140 658680 0 180 $X=830800 $Y=653260
X2397 4555 4562 2 1 4483 4557 MUX2 $T=835140 658680 1 180 $X=830800 $Y=658300
X2398 4567 4494 2 1 4546 4557 MUX2 $T=837620 688920 0 180 $X=833280 $Y=683500
X2399 4571 869 2 1 4598 4525 MUX2 $T=833900 578040 0 0 $X=833900 $Y=577660
X2400 4612 4609 2 1 4545 4537 MUX2 $T=840100 608280 1 180 $X=835760 $Y=607900
X2401 4603 869 2 1 4592 4625 MUX2 $T=838860 547800 0 0 $X=838860 $Y=547420
X2402 4632 4544 2 1 4547 871 MUX2 $T=843820 709080 1 180 $X=839480 $Y=708700
X2403 4622 879 2 1 4645 4525 MUX2 $T=841960 588120 1 0 $X=841960 $Y=582700
X2404 4636 869 2 1 4657 868 MUX2 $T=844440 567960 1 0 $X=844440 $Y=562540
X2405 4659 4658 2 1 4608 4537 MUX2 $T=848780 608280 1 180 $X=844440 $Y=607900
X2406 889 879 2 1 4614 4625 MUX2 $T=847540 547800 0 0 $X=847540 $Y=547420
X2407 4694 891 2 1 4726 4720 MUX2 $T=853740 567960 1 0 $X=853740 $Y=562540
X2408 4707 879 2 1 4735 4720 MUX2 $T=856220 578040 1 0 $X=856220 $Y=572620
X2409 4756 897 2 1 4775 4720 MUX2 $T=864280 567960 0 0 $X=864280 $Y=567580
X2410 4763 897 2 1 4785 4625 MUX2 $T=865520 557880 1 0 $X=865520 $Y=552460
X2411 4796 4731 2 1 4739 4760 MUX2 $T=871100 658680 0 180 $X=866760 $Y=653260
X2412 4773 914 2 1 4810 4759 MUX2 $T=868000 719160 0 0 $X=868000 $Y=718780
X2413 4811 4813 2 1 4784 4674 MUX2 $T=874820 598200 0 180 $X=870480 $Y=592780
X2414 4833 4731 2 1 4801 4767 MUX2 $T=879160 658680 0 180 $X=874820 $Y=653260
X2415 4815 4731 2 1 4823 4840 MUX2 $T=875440 628440 1 0 $X=875440 $Y=623020
X2416 4817 913 2 1 4841 4625 MUX2 $T=876060 547800 0 0 $X=876060 $Y=547420
X2417 4844 913 2 1 4781 922 MUX2 $T=881020 578040 1 180 $X=876680 $Y=577660
X2418 4824 913 2 1 4847 4720 MUX2 $T=877300 567960 0 0 $X=877300 $Y=567580
X2419 4779 4822 2 1 4866 4760 MUX2 $T=879780 648600 0 0 $X=879780 $Y=648220
X2420 927 4813 2 1 932 931 MUX2 $T=881640 537720 0 0 $X=881640 $Y=537340
X2421 4851 4813 2 1 4867 4625 MUX2 $T=881640 547800 0 0 $X=881640 $Y=547420
X2422 4854 4813 2 1 4876 4720 MUX2 $T=881640 567960 0 0 $X=881640 $Y=567580
X2423 4857 4813 2 1 4873 922 MUX2 $T=882260 578040 0 0 $X=882260 $Y=577660
X2424 4869 4822 2 1 4797 4767 MUX2 $T=884120 648600 0 0 $X=884120 $Y=648220
X2425 4909 4799 2 1 4864 816 MUX2 $T=890940 628440 0 180 $X=886600 $Y=623020
X2426 4919 4917 2 1 4838 4840 MUX2 $T=892800 547800 1 180 $X=888460 $Y=547420
X2427 4868 4701 2 1 4922 900 MUX2 $T=888460 688920 1 0 $X=888460 $Y=683500
X2428 4889 4943 2 1 4923 4767 MUX2 $T=897760 618360 1 180 $X=893420 $Y=617980
X2429 4879 4880 2 1 4911 4927 MUX2 $T=897760 688920 0 180 $X=893420 $Y=683500
X2430 4960 4888 2 1 4931 4515 MUX2 $T=900240 608280 0 180 $X=895900 $Y=602860
X2431 4964 4930 2 1 4937 821 MUX2 $T=901480 699000 1 180 $X=897140 $Y=698620
X2432 4978 4947 2 1 4938 4927 MUX2 $T=903960 648600 0 180 $X=899620 $Y=643180
X2433 958 4940 2 1 4941 807 MUX2 $T=904580 719160 1 180 $X=900240 $Y=718780
X2434 4961 4952 2 1 4985 4927 MUX2 $T=900860 688920 0 0 $X=900860 $Y=688540
X2435 4973 4955 2 1 4996 4949 MUX2 $T=902720 628440 0 0 $X=902720 $Y=628060
X2436 4995 4831 2 1 5027 4515 MUX2 $T=906440 598200 0 0 $X=906440 $Y=597820
X2437 5042 4925 2 1 4999 4966 MUX2 $T=913260 618360 0 180 $X=908920 $Y=612940
X2438 4828 4955 2 1 5006 4927 MUX2 $T=914500 638520 1 180 $X=910160 $Y=638140
X2439 5025 4957 2 1 5000 4927 MUX2 $T=914500 648600 1 180 $X=910160 $Y=648220
X2440 5028 4930 2 1 5052 968 MUX2 $T=910160 699000 0 0 $X=910160 $Y=698620
X2441 5029 4940 2 1 5049 968 MUX2 $T=910160 719160 1 0 $X=910160 $Y=713740
X2442 5056 4989 2 1 5048 4927 MUX2 $T=918220 668760 0 180 $X=913880 $Y=663340
X2443 5051 4947 2 1 5070 4949 MUX2 $T=914500 638520 0 0 $X=914500 $Y=638140
X2444 5061 4952 2 1 5072 4950 MUX2 $T=916360 688920 1 0 $X=916360 $Y=683500
X2445 5063 4957 2 1 5088 4949 MUX2 $T=916980 648600 0 0 $X=916980 $Y=648220
X2446 5081 4943 2 1 5067 4515 MUX2 $T=923180 598200 1 180 $X=918840 $Y=597820
X2447 979 4943 2 1 5077 4966 MUX2 $T=925040 608280 1 180 $X=920700 $Y=607900
X2448 5104 4940 2 1 5053 4759 MUX2 $T=925040 709080 0 180 $X=920700 $Y=703660
X2449 5076 4947 2 1 5126 5080 MUX2 $T=921320 648600 1 0 $X=921320 $Y=643180
X2450 5115 4989 2 1 5084 5080 MUX2 $T=926280 658680 1 180 $X=921940 $Y=658300
X2451 5096 4955 2 1 5141 5080 MUX2 $T=923800 628440 0 0 $X=923800 $Y=628060
X2452 5129 4930 2 1 5111 4759 MUX2 $T=930000 699000 1 180 $X=925660 $Y=698620
X2453 5033 4880 2 1 5085 4759 MUX2 $T=932480 678840 1 180 $X=928140 $Y=678460
X2454 5156 4989 2 1 5092 5131 MUX2 $T=933720 658680 0 180 $X=929380 $Y=653260
X2455 5147 4952 2 1 5176 5080 MUX2 $T=932480 678840 1 0 $X=932480 $Y=673420
X2456 5188 5151 2 1 5145 5155 MUX2 $T=939300 618360 0 180 $X=934960 $Y=612940
X2457 5189 4880 2 1 5135 992 MUX2 $T=939300 688920 0 180 $X=934960 $Y=683500
X2458 5143 4930 2 1 5185 992 MUX2 $T=935580 699000 0 0 $X=935580 $Y=698620
X2459 5180 4957 2 1 5204 5131 MUX2 $T=937440 658680 1 0 $X=937440 $Y=653260
X2460 5181 4957 2 1 5206 5080 MUX2 $T=938060 658680 0 0 $X=938060 $Y=658300
X2461 5190 4940 2 1 5197 992 MUX2 $T=938680 719160 1 0 $X=938680 $Y=713740
X2462 5198 4947 2 1 5223 5131 MUX2 $T=939920 638520 1 0 $X=939920 $Y=633100
X2463 5218 4952 2 1 5175 992 MUX2 $T=944260 678840 1 180 $X=939920 $Y=678460
X2464 5152 5151 2 1 5229 4966 MUX2 $T=941780 598200 0 0 $X=941780 $Y=597820
X2465 5210 4940 2 1 5241 936 MUX2 $T=943020 719160 1 0 $X=943020 $Y=713740
X2466 5236 5207 2 1 5257 4966 MUX2 $T=946120 598200 0 0 $X=946120 $Y=597820
X2467 5273 4930 2 1 5224 975 MUX2 $T=952320 699000 1 180 $X=947980 $Y=698620
X2468 5276 4877 2 1 5250 4966 MUX2 $T=952940 618360 0 180 $X=948600 $Y=612940
X2469 5256 4952 2 1 5281 5280 MUX2 $T=949220 688920 1 0 $X=949220 $Y=683500
X2470 1007 5284 2 1 5220 4966 MUX2 $T=954800 598200 1 180 $X=950460 $Y=597820
X2471 5262 4952 2 1 5286 5285 MUX2 $T=950460 678840 1 0 $X=950460 $Y=673420
X2472 5274 4940 2 1 5292 4423 MUX2 $T=952320 709080 1 0 $X=952320 $Y=703660
X2473 5279 4957 2 1 5294 5280 MUX2 $T=952940 658680 0 0 $X=952940 $Y=658300
X2474 5283 4957 2 1 5300 5285 MUX2 $T=954180 668760 1 0 $X=954180 $Y=663340
X2475 5287 4880 2 1 5301 5280 MUX2 $T=954180 688920 1 0 $X=954180 $Y=683500
X2476 5290 4955 2 1 5306 5285 MUX2 $T=956040 638520 0 0 $X=956040 $Y=638140
X2477 5291 4930 2 1 5309 4423 MUX2 $T=956040 699000 0 0 $X=956040 $Y=698620
X2478 5296 4877 2 1 5315 5312 MUX2 $T=957900 588120 1 0 $X=957900 $Y=582700
X2479 5317 5284 2 1 5298 4969 MUX2 $T=962240 618360 0 180 $X=957900 $Y=612940
X2480 5299 4989 2 1 5324 5280 MUX2 $T=957900 658680 0 0 $X=957900 $Y=658300
X2481 5304 4989 2 1 5322 5285 MUX2 $T=959140 668760 1 0 $X=959140 $Y=663340
X2482 5310 4947 2 1 5326 5280 MUX2 $T=961000 648600 1 0 $X=961000 $Y=643180
X2483 5320 5284 2 1 5333 5155 MUX2 $T=962860 608280 1 0 $X=962860 $Y=602860
X2484 5321 4877 2 1 5331 4969 MUX2 $T=962860 618360 1 0 $X=962860 $Y=612940
X2485 5325 5284 2 1 5340 5312 MUX2 $T=963480 588120 1 0 $X=963480 $Y=582700
X2486 5327 4880 2 1 5337 5285 MUX2 $T=964720 678840 1 0 $X=964720 $Y=673420
X2487 1022 4947 2 1 5323 5285 MUX2 $T=969680 648600 0 180 $X=965340 $Y=643180
X2488 5349 1024 2 1 5347 1029 MUX2 $T=972160 719160 0 0 $X=972160 $Y=718780
X2489 5365 4877 2 1 5382 5155 MUX2 $T=975260 598200 0 0 $X=975260 $Y=597820
X2490 5394 5368 2 1 5359 900 MUX2 $T=980840 699000 0 180 $X=976500 $Y=693580
X2491 5401 5350 2 1 5351 4969 MUX2 $T=981460 638520 0 180 $X=977120 $Y=633100
X2492 5355 5345 2 1 5332 5312 MUX2 $T=983320 588120 1 180 $X=978980 $Y=587740
X2493 5361 5420 2 1 5399 1034 MUX2 $T=986420 598200 1 180 $X=982080 $Y=597820
X2494 5430 5350 2 1 5405 816 MUX2 $T=987040 638520 0 180 $X=982700 $Y=633100
X2495 5416 5412 2 1 5452 4969 MUX2 $T=984560 618360 0 0 $X=984560 $Y=617980
X2496 1063 5467 2 1 5484 5458 MUX2 $T=991380 567960 0 0 $X=991380 $Y=567580
X2497 5486 5420 2 1 5363 5445 MUX2 $T=995720 608280 1 180 $X=991380 $Y=607900
X2498 5465 5466 2 1 5489 5477 MUX2 $T=992000 648600 0 0 $X=992000 $Y=648220
X2499 5503 5469 2 1 5418 5477 MUX2 $T=997580 678840 1 180 $X=993240 $Y=678460
X2500 5569 5522 2 1 5546 5445 MUX2 $T=1009360 608280 0 180 $X=1005020 $Y=602860
X2501 5622 5547 2 1 5644 5445 MUX2 $T=1016180 588120 0 0 $X=1016180 $Y=587740
X2502 5658 5420 2 1 5606 5155 MUX2 $T=1022380 608280 1 180 $X=1018040 $Y=607900
X2503 5651 5654 2 1 5661 5650 MUX2 $T=1021760 608280 1 0 $X=1021760 $Y=602860
X2504 5675 5619 2 1 5694 1097 MUX2 $T=1026100 578040 1 0 $X=1026100 $Y=572620
X2505 5703 5522 2 1 5670 5650 MUX2 $T=1031060 608280 0 180 $X=1026720 $Y=602860
X2506 5691 5638 2 1 5695 1097 MUX2 $T=1034780 578040 0 180 $X=1030440 $Y=572620
X2507 5752 5494 2 1 5726 5650 MUX2 $T=1042220 608280 1 180 $X=1037880 $Y=607900
X2508 5783 5778 2 1 5758 5760 MUX2 $T=1047180 578040 1 180 $X=1042840 $Y=577660
X2509 5767 5610 2 1 5787 5781 MUX2 $T=1043460 699000 0 0 $X=1043460 $Y=698620
X2510 5769 5763 2 1 5772 5760 MUX2 $T=1049040 567960 1 180 $X=1044700 $Y=567580
X2511 5776 5612 2 1 5798 5797 MUX2 $T=1045320 658680 1 0 $X=1045320 $Y=653260
X2512 5779 5774 2 1 5799 1123 MUX2 $T=1045940 608280 0 0 $X=1045940 $Y=607900
X2513 5786 5771 2 1 5804 5797 MUX2 $T=1047180 628440 0 0 $X=1047180 $Y=628060
X2514 5807 5443 2 1 5788 5760 MUX2 $T=1052140 567960 0 180 $X=1047800 $Y=562540
X2515 5789 5625 2 1 5727 5797 MUX2 $T=1047800 618360 0 0 $X=1047800 $Y=617980
X2516 5793 5448 2 1 1126 1129 MUX2 $T=1049040 537720 0 0 $X=1049040 $Y=537340
X2517 5816 5782 2 1 5795 1123 MUX2 $T=1053380 598200 0 180 $X=1049040 $Y=592780
X2518 5844 5751 2 1 5819 1127 MUX2 $T=1057720 588120 1 180 $X=1053380 $Y=587740
X2519 5850 5842 2 1 5815 1128 MUX2 $T=1058340 547800 1 180 $X=1054000 $Y=547420
X2520 5851 5826 2 1 5831 1123 MUX2 $T=1058960 598200 0 180 $X=1054620 $Y=592780
X2521 5832 5813 2 1 5854 5858 MUX2 $T=1054620 699000 1 0 $X=1054620 $Y=693580
X2522 5835 1130 2 1 5834 1118 MUX2 $T=1058960 719160 1 180 $X=1054620 $Y=718780
X2523 5860 5838 2 1 5805 5732 MUX2 $T=1059580 628440 1 180 $X=1055240 $Y=628060
X2524 5862 5751 2 1 5821 5797 MUX2 $T=1061440 608280 1 180 $X=1057100 $Y=607900
X2525 5796 5845 2 1 5802 5732 MUX2 $T=1061440 648600 1 180 $X=1057100 $Y=648220
X2526 5666 5842 2 1 5870 1133 MUX2 $T=1058960 547800 1 0 $X=1058960 $Y=542380
X2527 1131 5778 2 1 5888 1133 MUX2 $T=1058960 547800 0 0 $X=1058960 $Y=547420
X2528 5873 5812 2 1 5808 5732 MUX2 $T=1063300 668760 0 180 $X=1058960 $Y=663340
X2529 5901 5887 2 1 5809 5732 MUX2 $T=1067640 678840 0 180 $X=1063300 $Y=673420
X2530 1137 1134 2 1 5907 1142 MUX2 $T=1065780 719160 0 0 $X=1065780 $Y=718780
X2531 5913 5774 2 1 5881 4949 MUX2 $T=1070740 618360 0 180 $X=1066400 $Y=612940
X2532 5895 5826 2 1 5830 1127 MUX2 $T=1067020 578040 0 0 $X=1067020 $Y=577660
X2533 5875 5794 2 1 5917 1133 MUX2 $T=1067640 557880 0 0 $X=1067640 $Y=557500
X2534 5876 5845 2 1 5920 5897 MUX2 $T=1067640 658680 1 0 $X=1067640 $Y=653260
X2535 5903 5782 2 1 5919 1127 MUX2 $T=1068260 598200 0 0 $X=1068260 $Y=597820
X2536 5892 5751 2 1 5926 1140 MUX2 $T=1069500 588120 1 0 $X=1069500 $Y=582700
X2537 5915 5813 2 1 5918 5890 MUX2 $T=1071360 699000 0 0 $X=1071360 $Y=698620
X2538 5930 5806 2 1 5947 5890 MUX2 $T=1073220 709080 1 0 $X=1073220 $Y=703660
X2539 1150 5842 2 1 5934 1146 MUX2 $T=1078800 547800 0 180 $X=1074460 $Y=542380
X2540 5952 5853 2 1 5905 5890 MUX2 $T=1078800 678840 1 180 $X=1074460 $Y=678460
X2541 5931 5778 2 1 5954 1140 MUX2 $T=1075080 557880 0 0 $X=1075080 $Y=557500
X2542 5958 5774 2 1 5942 1146 MUX2 $T=1080660 608280 1 180 $X=1076320 $Y=607900
X2543 5965 5806 2 1 5950 1142 MUX2 $T=1081900 709080 0 180 $X=1077560 $Y=703660
X2544 1154 5763 2 1 5955 1140 MUX2 $T=1083140 567960 1 180 $X=1078800 $Y=567580
X2545 5971 5853 2 1 5941 5946 MUX2 $T=1083140 658680 1 180 $X=1078800 $Y=658300
X2546 5959 5853 2 1 5984 1156 MUX2 $T=1080660 688920 0 0 $X=1080660 $Y=688540
X2547 5980 5771 2 1 5948 5946 MUX2 $T=1085620 628440 1 180 $X=1081280 $Y=628060
X2548 5997 5845 2 1 5967 1156 MUX2 $T=1088100 678840 0 180 $X=1083760 $Y=673420
X2549 5985 5794 2 1 6004 1140 MUX2 $T=1085620 557880 1 0 $X=1085620 $Y=552460
X2550 5987 5853 2 1 5983 1142 MUX2 $T=1085620 668760 1 0 $X=1085620 $Y=663340
X2551 6031 5782 2 1 5972 5995 MUX2 $T=1091820 608280 0 180 $X=1087480 $Y=602860
X2552 5966 5845 2 1 6018 5946 MUX2 $T=1087480 648600 0 0 $X=1087480 $Y=648220
X2553 6011 5806 2 1 6048 6013 MUX2 $T=1090580 699000 1 0 $X=1090580 $Y=693580
X2554 6010 5838 2 1 6033 6005 MUX2 $T=1091200 628440 1 0 $X=1091200 $Y=623020
X2555 6020 5794 2 1 5964 5995 MUX2 $T=1092440 557880 1 0 $X=1092440 $Y=552460
X2556 6026 5845 2 1 6063 6005 MUX2 $T=1093060 648600 0 0 $X=1093060 $Y=648220
X2557 6006 5838 2 1 6059 6056 MUX2 $T=1093680 618360 1 0 $X=1093680 $Y=612940
X2558 6035 5782 2 1 6040 6056 MUX2 $T=1094300 588120 1 0 $X=1094300 $Y=582700
X2559 6039 5771 2 1 6087 6005 MUX2 $T=1095540 628440 1 0 $X=1095540 $Y=623020
X2560 6052 1134 2 1 6084 1156 MUX2 $T=1096780 719160 0 0 $X=1096780 $Y=718780
X2561 1170 5842 2 1 6076 6075 MUX2 $T=1098020 547800 1 0 $X=1098020 $Y=542380
X2562 6083 5813 2 1 6036 1142 MUX2 $T=1102360 699000 1 180 $X=1098020 $Y=698620
X2563 6060 5774 2 1 6081 6056 MUX2 $T=1098640 588120 1 0 $X=1098640 $Y=582700
X2564 6065 5774 2 1 6093 5995 MUX2 $T=1099880 618360 1 0 $X=1099880 $Y=612940
X2565 6099 5887 2 1 6046 6077 MUX2 $T=1106080 668760 1 180 $X=1101740 $Y=668380
X2566 1174 5842 2 1 6102 6101 MUX2 $T=1102360 547800 1 0 $X=1102360 $Y=542380
X2567 6112 5812 2 1 6086 6013 MUX2 $T=1107320 668760 0 180 $X=1102980 $Y=663340
X2568 6115 5887 2 1 6088 6013 MUX2 $T=1107940 658680 1 180 $X=1103600 $Y=658300
X2569 6116 5813 2 1 6095 6013 MUX2 $T=1107940 699000 0 180 $X=1103600 $Y=693580
X2570 6097 5838 2 1 6123 6013 MUX2 $T=1105460 638520 1 0 $X=1105460 $Y=633100
X2571 6078 1134 2 1 6124 1135 MUX2 $T=1105460 719160 0 0 $X=1105460 $Y=718780
X2572 6109 5794 2 1 6130 6075 MUX2 $T=1106700 547800 1 0 $X=1106700 $Y=542380
X2573 6120 5813 2 1 6144 1183 MUX2 $T=1107940 699000 1 0 $X=1107940 $Y=693580
X2574 6121 5763 2 1 6165 6138 MUX2 $T=1108560 618360 1 0 $X=1108560 $Y=612940
X2575 1182 5763 2 1 6152 6075 MUX2 $T=1109180 567960 0 0 $X=1109180 $Y=567580
X2576 6126 5778 2 1 6169 6138 MUX2 $T=1110420 598200 0 0 $X=1110420 $Y=597820
X2577 6127 5751 2 1 6161 6138 MUX2 $T=1110420 608280 1 0 $X=1110420 $Y=602860
X2578 6132 5771 2 1 6155 6013 MUX2 $T=1110420 638520 1 0 $X=1110420 $Y=633100
X2579 6134 1134 2 1 6162 1183 MUX2 $T=1110420 719160 0 0 $X=1110420 $Y=718780
X2580 6136 5826 2 1 6154 6056 MUX2 $T=1111040 588120 1 0 $X=1111040 $Y=582700
X2581 6137 5826 2 1 6157 6101 MUX2 $T=1111040 598200 1 0 $X=1111040 $Y=592780
X2582 6085 5778 2 1 6166 6101 MUX2 $T=1112280 567960 1 0 $X=1112280 $Y=562540
X2583 6147 5826 2 1 6176 6138 MUX2 $T=1112280 608280 0 0 $X=1112280 $Y=607900
X2584 6148 5812 2 1 6167 6077 MUX2 $T=1112280 668760 1 0 $X=1112280 $Y=663340
X2585 6150 5887 2 1 6047 6140 MUX2 $T=1112280 678840 0 0 $X=1112280 $Y=678460
X2586 6151 5806 2 1 6171 1183 MUX2 $T=1112280 699000 1 0 $X=1112280 $Y=693580
X2587 6145 5806 2 1 6168 6140 MUX2 $T=1112280 699000 0 0 $X=1112280 $Y=698620
X2588 6096 5887 2 1 6170 5946 MUX2 $T=1112900 658680 1 0 $X=1112900 $Y=653260
X2589 6153 5763 2 1 6172 6101 MUX2 $T=1114140 567960 0 0 $X=1114140 $Y=567580
X2590 6156 5812 2 1 6175 6140 MUX2 $T=1114140 678840 1 0 $X=1114140 $Y=673420
X2591 6158 5771 2 1 6177 6140 MUX2 $T=1114760 638520 1 0 $X=1114760 $Y=633100
X2592 6163 5751 2 1 6173 6101 MUX2 $T=1115380 588120 1 0 $X=1115380 $Y=582700
X2593 6174 5812 2 1 6180 5946 MUX2 $T=1117860 658680 1 0 $X=1117860 $Y=653260
X2594 6179 5778 2 1 6183 6075 MUX2 $T=1121580 557880 1 0 $X=1121580 $Y=552460
X2595 1804 1762 1776 1796 1 1772 2 AOI22S $T=322400 598200 0 0 $X=322400 $Y=597820
X2596 2051 2040 1951 2009 1 2018 2 AOI22S $T=372620 688920 0 180 $X=368900 $Y=683500
X2597 2051 2031 191 2009 1 2058 2 AOI22S $T=372000 678840 1 0 $X=372000 $Y=673420
X2598 2051 2026 192 2009 1 2045 2 AOI22S $T=376340 688920 0 180 $X=372620 $Y=683500
X2599 2051 2093 2096 2009 1 1991 2 AOI22S $T=381920 688920 0 180 $X=378200 $Y=683500
X2600 2051 2061 203 2116 1 2107 2 AOI22S $T=386880 668760 0 180 $X=383160 $Y=663340
X2601 2051 2124 2121 2009 1 2131 2 AOI22S $T=384400 678840 0 0 $X=384400 $Y=678460
X2602 2139 2142 212 2116 1 2194 2 AOI22S $T=401140 668760 0 180 $X=397420 $Y=663340
X2603 2139 2198 213 2116 1 2179 2 AOI22S $T=400520 668760 0 0 $X=400520 $Y=668380
X2604 2116 2226 2227 2139 1 2186 2 AOI22S $T=404860 668760 0 180 $X=401140 $Y=663340
X2605 2116 2273 222 2139 1 2252 2 AOI22S $T=412920 668760 0 0 $X=412920 $Y=668380
X2606 2322 2306 2317 2301 1 2129 2 AOI22S $T=420980 648600 1 180 $X=417260 $Y=648220
X2607 2322 2330 2342 2301 1 2173 2 AOI22S $T=424700 658680 0 180 $X=420980 $Y=653260
X2608 2322 2255 2366 2301 1 2135 2 AOI22S $T=428420 658680 0 180 $X=424700 $Y=653260
X2609 2401 2314 2391 2387 1 2305 2 AOI22S $T=432760 648600 0 180 $X=429040 $Y=643180
X2610 2322 2402 245 2301 1 2243 2 AOI22S $T=435240 658680 0 180 $X=431520 $Y=653260
X2611 2322 2442 253 2301 1 2219 2 AOI22S $T=442060 658680 1 180 $X=438340 $Y=658300
X2612 2401 2484 2485 2387 1 2388 2 AOI22S $T=448880 648600 0 180 $X=445160 $Y=643180
X2613 2322 2487 256 2481 1 2356 2 AOI22S $T=446400 648600 0 0 $X=446400 $Y=648220
X2614 2474 2518 2516 2504 1 2413 2 AOI22S $T=452600 648600 1 0 $X=452600 $Y=643180
X2615 2401 2561 2544 2481 1 2389 2 AOI22S $T=458800 648600 1 0 $X=458800 $Y=643180
X2616 2547 2586 2597 2539 1 2172 2 AOI22S $T=466240 608280 0 180 $X=462520 $Y=602860
X2617 2868 2858 359 2811 1 2818 2 AOI22S $T=515220 719160 0 180 $X=511500 $Y=713740
X2618 2868 2858 362 2874 1 2795 2 AOI22S $T=515220 709080 0 0 $X=515220 $Y=708700
X2619 2889 2858 367 2886 1 371 2 AOI22S $T=519560 719160 0 0 $X=519560 $Y=718780
X2620 2889 2962 386 2965 1 2934 2 AOI22S $T=530100 709080 0 0 $X=530100 $Y=708700
X2621 2889 2962 419 409 1 412 2 AOI22S $T=554280 719160 0 180 $X=550560 $Y=713740
X2622 2889 2962 422 3059 1 3093 2 AOI22S $T=553660 709080 0 0 $X=553660 $Y=708700
X2623 433 2962 446 2681 1 2949 2 AOI22S $T=563580 709080 0 0 $X=563580 $Y=708700
X2624 433 452 469 466 1 3178 2 AOI22S $T=572260 719160 1 0 $X=572260 $Y=713740
X2625 433 452 486 3204 1 491 2 AOI22S $T=581560 719160 1 0 $X=581560 $Y=713740
X2626 580 573 577 538 1 2931 2 AOI22S $T=616900 719160 1 180 $X=613180 $Y=718780
X2627 3452 3423 3422 3421 1 3436 2 AOI22S $T=624960 688920 1 180 $X=621240 $Y=688540
X2628 580 573 623 621 1 2885 2 AOI22S $T=641080 719160 0 180 $X=637360 $Y=713740
X2629 3615 3607 3619 3577 1 3526 2 AOI22S $T=652860 658680 1 180 $X=649140 $Y=658300
X2630 3615 3607 3617 3589 1 3565 2 AOI22S $T=653480 618360 0 180 $X=649760 $Y=612940
X2631 3615 3607 3618 3558 1 3402 2 AOI22S $T=653480 648600 1 180 $X=649760 $Y=648220
X2632 3615 3607 3638 3631 1 3121 2 AOI22S $T=657820 658680 1 180 $X=654100 $Y=658300
X2633 3660 3607 3651 3559 1 3586 2 AOI22S $T=660300 668760 1 180 $X=656580 $Y=668380
X2634 3615 3654 3675 3569 1 3266 2 AOI22S $T=662780 608280 0 180 $X=659060 $Y=602860
X2635 3681 3654 3674 3614 1 3616 2 AOI22S $T=663400 598200 1 180 $X=659680 $Y=597820
X2636 3660 3607 3688 3666 1 3662 2 AOI22S $T=663400 678840 1 180 $X=659680 $Y=678460
X2637 3681 3654 3673 3649 1 3622 2 AOI22S $T=664020 588120 0 180 $X=660300 $Y=582700
X2638 3681 661 665 662 1 3691 2 AOI22S $T=672700 537720 1 180 $X=668980 $Y=537340
X2639 3681 661 3745 3449 1 3698 2 AOI22S $T=672700 567960 0 180 $X=668980 $Y=562540
X2640 3742 3723 3729 3682 1 3611 2 AOI22S $T=672700 638520 1 180 $X=668980 $Y=638140
X2641 3730 3725 3734 3696 1 3643 2 AOI22S $T=672700 668760 1 180 $X=668980 $Y=668380
X2642 3742 3723 3758 3420 1 3647 2 AOI22S $T=677040 638520 1 180 $X=673320 $Y=638140
X2643 3771 3760 3737 3719 1 3753 2 AOI22S $T=679520 688920 1 180 $X=675800 $Y=688540
X2644 3788 3774 3782 3703 1 3773 2 AOI22S $T=682620 608280 0 180 $X=678900 $Y=602860
X2645 3788 3774 3784 3770 1 3735 2 AOI22S $T=683240 598200 0 180 $X=679520 $Y=592780
X2646 681 3786 3789 3336 1 3780 2 AOI22S $T=684480 567960 0 180 $X=680760 $Y=562540
X2647 681 680 3794 3762 1 3393 2 AOI22S $T=685720 557880 0 180 $X=682000 $Y=552460
X2648 3742 3723 3795 3748 1 3582 2 AOI22S $T=685720 638520 1 180 $X=682000 $Y=638140
X2649 3730 3725 3808 3790 1 3041 2 AOI22S $T=686340 658680 1 180 $X=682620 $Y=658300
X2650 3730 3725 3801 3796 1 3777 2 AOI22S $T=686960 668760 1 180 $X=683240 $Y=668380
X2651 681 680 3817 673 1 3598 2 AOI22S $T=690060 557880 0 180 $X=686340 $Y=552460
X2652 3820 3786 3802 3599 1 3492 2 AOI22S $T=690060 588120 0 180 $X=686340 $Y=582700
X2653 3788 3774 3818 3194 1 3672 2 AOI22S $T=690060 598200 1 180 $X=686340 $Y=597820
X2654 639 687 689 686 1 3809 2 AOI22S $T=690060 719160 1 180 $X=686340 $Y=718780
X2655 3771 3760 3812 3112 1 3805 2 AOI22S $T=687580 688920 0 0 $X=687580 $Y=688540
X2656 3771 3760 3810 3837 1 3294 2 AOI22S $T=691300 688920 0 0 $X=691300 $Y=688540
X2657 3742 3723 3857 3793 1 3827 2 AOI22S $T=696260 638520 1 180 $X=692540 $Y=638140
X2658 3855 3859 3830 3671 1 3787 2 AOI22S $T=698120 567960 1 180 $X=694400 $Y=567580
X2659 3788 3774 3869 3850 1 3821 2 AOI22S $T=698120 598200 1 180 $X=694400 $Y=597820
X2660 3730 3725 3852 3815 1 3886 2 AOI22S $T=698120 668760 1 0 $X=698120 $Y=663340
X2661 699 702 3835 3881 1 3653 2 AOI22S $T=698740 557880 1 0 $X=698740 $Y=552460
X2662 3788 3774 3895 3552 1 3286 2 AOI22S $T=703700 608280 1 0 $X=703700 $Y=602860
X2663 3855 3903 3899 3447 1 3887 2 AOI22S $T=705560 567960 0 0 $X=705560 $Y=567580
X2664 3820 3786 3908 3904 1 3686 2 AOI22S $T=710520 588120 1 180 $X=706800 $Y=587740
X2665 3730 3725 3910 3898 1 3208 2 AOI22S $T=710520 668760 1 180 $X=706800 $Y=668380
X2666 3873 3859 3919 3907 1 3625 2 AOI22S $T=712380 638520 1 180 $X=708660 $Y=638140
X2667 3771 3760 3915 3102 1 3018 2 AOI22S $T=709900 688920 1 0 $X=709900 $Y=683500
X2668 3730 3725 3981 3868 1 3917 2 AOI22S $T=722300 668760 1 180 $X=718580 $Y=668380
X2669 3855 3903 3921 3970 1 3945 2 AOI22S $T=720440 557880 1 0 $X=720440 $Y=552460
X2670 3660 3979 3982 3963 1 3969 2 AOI22S $T=724160 678840 0 180 $X=720440 $Y=673420
X2671 705 708 3987 3950 1 3938 2 AOI22S $T=724780 608280 1 180 $X=721060 $Y=607900
X2672 3820 3786 3977 3956 1 3924 2 AOI22S $T=723540 588120 0 0 $X=723540 $Y=587740
X2673 3873 3859 4004 3933 1 3993 2 AOI22S $T=727880 638520 1 180 $X=724160 $Y=638140
X2674 3771 3760 3994 3999 1 4000 2 AOI22S $T=724160 688920 0 0 $X=724160 $Y=688540
X2675 3992 3728 3991 3973 1 4003 2 AOI22S $T=724780 618360 1 0 $X=724780 $Y=612940
X2676 4019 3996 4081 4036 1 3301 2 AOI22S $T=740900 648600 1 180 $X=737180 $Y=648220
X2677 3820 3786 4088 4063 1 3906 2 AOI22S $T=742140 598200 0 180 $X=738420 $Y=592780
X2678 4080 3978 4098 3990 1 4001 2 AOI22S $T=746480 668760 1 180 $X=742760 $Y=668380
X2679 3992 3728 4146 4128 1 4136 2 AOI22S $T=756400 608280 1 180 $X=752680 $Y=607900
X2680 4025 708 4147 3154 1 4137 2 AOI22S $T=756400 628440 0 180 $X=752680 $Y=623020
X2681 4134 774 4151 4092 1 3515 2 AOI22S $T=757020 567960 1 180 $X=753300 $Y=567580
X2682 4134 774 4154 4142 1 4085 2 AOI22S $T=757640 547800 1 180 $X=753920 $Y=547420
X2683 4134 774 4161 3341 1 4045 2 AOI22S $T=757640 557880 1 180 $X=753920 $Y=557500
X2684 4080 3996 4163 4119 1 3483 2 AOI22S $T=758260 658680 1 180 $X=754540 $Y=658300
X2685 3820 774 4152 4141 1 3455 2 AOI22S $T=755160 588120 0 0 $X=755160 $Y=587740
X2686 4080 3978 4166 4158 1 4139 2 AOI22S $T=758880 668760 1 180 $X=755160 $Y=668380
X2687 4080 3996 4186 3378 1 4162 2 AOI22S $T=760120 648600 0 180 $X=756400 $Y=643180
X2688 4080 3978 4189 4130 1 3259 2 AOI22S $T=760740 658680 0 0 $X=760740 $Y=658300
X2689 4218 4180 4206 4199 1 4160 2 AOI22S $T=767560 688920 0 180 $X=763840 $Y=683500
X2690 3992 3728 4215 4191 1 4179 2 AOI22S $T=768800 598200 1 180 $X=765080 $Y=597820
X2691 3992 3979 4224 4214 1 4213 2 AOI22S $T=770040 578040 1 180 $X=766320 $Y=577660
X2692 4208 4216 4202 3560 1 4226 2 AOI22S $T=766320 699000 0 0 $X=766320 $Y=698620
X2693 4025 4106 4231 4093 1 4086 2 AOI22S $T=771280 608280 0 0 $X=771280 $Y=607900
X2694 801 798 799 797 1 751 2 AOI22S $T=776860 537720 1 180 $X=773140 $Y=537340
X2695 3660 4260 4263 4256 1 3451 2 AOI22S $T=778100 668760 1 180 $X=774380 $Y=668380
X2696 4208 4216 4272 4234 1 4255 2 AOI22S $T=779340 699000 1 180 $X=775620 $Y=698620
X2697 808 793 4302 4270 1 4257 2 AOI22S $T=783680 547800 1 180 $X=779960 $Y=547420
X2698 4258 4254 4241 4277 1 4264 2 AOI22S $T=779960 598200 0 0 $X=779960 $Y=597820
X2699 4283 4294 4286 4296 1 4300 2 AOI22S $T=781200 648600 0 0 $X=781200 $Y=648220
X2700 808 793 4303 4295 1 3496 2 AOI22S $T=785540 557880 1 180 $X=781820 $Y=557500
X2701 4025 4106 4267 4291 1 4127 2 AOI22S $T=781820 618360 1 0 $X=781820 $Y=612940
X2702 3992 793 4306 3639 1 4250 2 AOI22S $T=786160 588120 0 180 $X=782440 $Y=582700
X2703 4218 4260 4314 4301 1 3293 2 AOI22S $T=789880 678840 0 180 $X=786160 $Y=673420
X2704 4208 4216 4309 4284 1 3298 2 AOI22S $T=786160 699000 1 0 $X=786160 $Y=693580
X2705 4258 4254 4276 3476 1 4280 2 AOI22S $T=791740 578040 0 180 $X=788020 $Y=572620
X2706 4258 4254 4311 4337 1 4334 2 AOI22S $T=792980 588120 0 180 $X=789260 $Y=582700
X2707 801 4106 4298 3522 1 4344 2 AOI22S $T=789880 598200 0 0 $X=789880 $Y=597820
X2708 4218 4260 4346 3323 1 3389 2 AOI22S $T=793600 678840 1 180 $X=789880 $Y=678460
X2709 4208 4216 4336 3281 1 4352 2 AOI22S $T=791120 699000 1 0 $X=791120 $Y=693580
X2710 4258 4254 4312 4355 1 4351 2 AOI22S $T=793600 598200 1 0 $X=793600 $Y=592780
X2711 4258 4254 4363 4371 1 4319 2 AOI22S $T=796080 567960 1 0 $X=796080 $Y=562540
X2712 4208 4216 4364 4375 1 3344 2 AOI22S $T=796080 699000 1 0 $X=796080 $Y=693580
X2713 4283 4294 4368 3462 1 4382 2 AOI22S $T=796700 648600 1 0 $X=796700 $Y=643180
X2714 4218 4260 4369 4379 1 3370 2 AOI22S $T=796700 678840 1 0 $X=796700 $Y=673420
X2715 4218 4260 4374 4383 1 3435 2 AOI22S $T=797320 678840 0 0 $X=797320 $Y=678460
X2716 4283 4294 4391 3327 1 4361 2 AOI22S $T=800420 648600 0 0 $X=800420 $Y=648220
X2717 4208 4216 4392 3443 1 4399 2 AOI22S $T=800420 699000 0 0 $X=800420 $Y=698620
X2718 801 798 825 4376 1 826 2 AOI22S $T=802900 537720 0 0 $X=802900 $Y=537340
X2719 4534 4523 4527 4517 1 4462 2 AOI22S $T=828320 699000 0 180 $X=824600 $Y=693580
X2720 4566 4561 4516 3433 1 3461 2 AOI22S $T=833280 668760 1 180 $X=829560 $Y=668380
X2721 870 866 4597 4559 1 4425 2 AOI22S $T=835760 547800 1 180 $X=832040 $Y=547420
X2722 4591 4573 4533 4538 1 4502 2 AOI22S $T=836380 638520 1 180 $X=832660 $Y=638140
X2723 870 4577 4584 4569 1 4560 2 AOI22S $T=837000 588120 0 180 $X=833280 $Y=582700
X2724 870 866 4587 4496 1 4512 2 AOI22S $T=837620 567960 1 180 $X=833900 $Y=567580
X2725 4591 4588 4596 3523 1 4539 2 AOI22S $T=838240 648600 1 180 $X=834520 $Y=648220
X2726 4534 4523 4593 4491 1 4581 2 AOI22S $T=838240 699000 0 180 $X=834520 $Y=693580
X2727 4583 4588 4602 4520 1 4549 2 AOI22S $T=839480 658680 1 180 $X=835760 $Y=658300
X2728 4534 4604 4600 4575 1 4506 2 AOI22S $T=837620 608280 1 0 $X=837620 $Y=602860
X2729 4591 4588 4616 4536 1 4606 2 AOI22S $T=841960 578040 1 180 $X=838240 $Y=577660
X2730 4591 4573 4629 875 1 3547 2 AOI22S $T=843820 638520 1 180 $X=840100 $Y=638140
X2731 4591 4573 4628 4621 1 4619 2 AOI22S $T=844440 608280 1 180 $X=840720 $Y=607900
X2732 886 885 4646 4518 1 865 2 AOI22S $T=847540 547800 1 180 $X=843820 $Y=547420
X2733 4566 4561 4641 4509 1 4624 2 AOI22S $T=845680 668760 0 0 $X=845680 $Y=668380
X2734 4534 4523 4648 4656 1 4664 2 AOI22S $T=846300 699000 1 0 $X=846300 $Y=693580
X2735 886 885 4667 4613 1 4677 2 AOI22S $T=849400 567960 1 0 $X=849400 $Y=562540
X2736 4583 4588 4698 4670 1 4686 2 AOI22S $T=856220 658680 0 180 $X=852500 $Y=653260
X2737 4679 4692 4700 4693 1 4691 2 AOI22S $T=856220 699000 0 180 $X=852500 $Y=693580
X2738 4690 4703 4721 4709 1 4716 2 AOI22S $T=856840 678840 1 0 $X=856840 $Y=673420
X2739 4708 4718 4618 4711 1 4678 2 AOI22S $T=857460 588120 0 0 $X=857460 $Y=587740
X2740 4708 901 4680 4734 1 4696 2 AOI22S $T=863660 567960 1 180 $X=859940 $Y=567580
X2741 4477 4743 4510 4688 1 4728 2 AOI22S $T=863660 648600 0 180 $X=859940 $Y=643180
X2742 4757 4743 4729 4736 1 4697 2 AOI22S $T=866140 648600 1 180 $X=862420 $Y=648220
X2743 4679 4692 4750 4755 1 4762 2 AOI22S $T=862420 699000 1 0 $X=862420 $Y=693580
X2744 4757 4743 4586 4782 1 4780 2 AOI22S $T=866140 648600 0 0 $X=866140 $Y=648220
X2745 917 919 4644 4787 1 4798 2 AOI22S $T=869860 557880 1 0 $X=869860 $Y=552460
X2746 4690 4703 4771 4793 1 4791 2 AOI22S $T=869860 678840 1 0 $X=869860 $Y=673420
X2747 917 4500 4687 4794 1 4800 2 AOI22S $T=870480 567960 0 0 $X=870480 $Y=567580
X2748 4477 4500 4649 4774 1 4808 2 AOI22S $T=871720 598200 0 0 $X=871720 $Y=597820
X2749 917 4500 4611 4806 1 4807 2 AOI22S $T=872340 578040 0 0 $X=872340 $Y=577660
X2750 4795 4803 4777 4764 1 4790 2 AOI22S $T=872340 648600 0 0 $X=872340 $Y=648220
X2751 4795 4803 4843 4845 1 4859 2 AOI22S $T=879780 658680 1 0 $X=879780 $Y=653260
X2752 4679 4692 4861 4846 1 4858 2 AOI22S $T=885360 699000 0 180 $X=881640 $Y=693580
X2753 4583 4573 4872 4885 1 4882 2 AOI22S $T=884740 658680 0 0 $X=884740 $Y=658300
X2754 4690 4703 4853 4834 1 4893 2 AOI22S $T=885360 668760 0 0 $X=885360 $Y=668380
X2755 4915 4905 4908 4829 1 4899 2 AOI22S $T=891560 608280 1 180 $X=887840 $Y=607900
X2756 4915 4905 4934 4821 1 4914 2 AOI22S $T=895900 608280 0 180 $X=892180 $Y=602860
X2757 4915 4905 4975 4953 1 4956 2 AOI22S $T=904580 608280 0 180 $X=900860 $Y=602860
X2758 4990 4976 4982 944 1 953 2 AOI22S $T=905200 557880 0 180 $X=901480 $Y=552460
X2759 4679 4692 4980 4971 1 952 2 AOI22S $T=905200 699000 1 180 $X=901480 $Y=698620
X2760 4915 4905 4994 955 1 4954 2 AOI22S $T=905820 567960 0 180 $X=902100 $Y=562540
X2761 4795 4884 4965 4802 1 4987 2 AOI22S $T=902720 638520 0 0 $X=902720 $Y=638140
X2762 4690 4703 4981 4842 1 4951 2 AOI22S $T=907680 688920 0 180 $X=903960 $Y=683500
X2763 4915 4905 4992 948 1 5009 2 AOI22S $T=905200 578040 0 0 $X=905200 $Y=577660
X2764 4912 4998 5005 4920 1 4862 2 AOI22S $T=908920 618360 0 180 $X=905200 $Y=612940
X2765 4679 4692 4988 5013 1 5004 2 AOI22S $T=905820 699000 0 0 $X=905820 $Y=698620
X2766 4795 4884 4970 5014 1 5015 2 AOI22S $T=906440 638520 0 0 $X=906440 $Y=638140
X2767 4990 4976 5019 959 1 4916 2 AOI22S $T=910780 547800 1 180 $X=907060 $Y=547420
X2768 4963 5021 4997 5018 1 5034 2 AOI22S $T=909540 668760 1 0 $X=909540 $Y=663340
X2769 5071 4786 5064 5001 1 967 2 AOI22S $T=918840 547800 1 180 $X=915120 $Y=547420
X2770 4912 4998 5065 5068 1 971 2 AOI22S $T=916980 618360 1 0 $X=916980 $Y=612940
X2771 5071 4786 5074 5008 1 973 2 AOI22S $T=918840 547800 0 0 $X=918840 $Y=547420
X2772 4912 4786 5083 5046 1 5038 2 AOI22S $T=923180 567960 0 180 $X=919460 $Y=562540
X2773 4912 4786 5086 5058 1 5095 2 AOI22S $T=921320 588120 1 0 $X=921320 $Y=582700
X2774 5007 5103 5093 5098 1 5110 2 AOI22S $T=923180 699000 1 0 $X=923180 $Y=693580
X2775 5102 5089 5106 5003 1 5116 2 AOI22S $T=924420 678840 0 0 $X=924420 $Y=678460
X2776 5091 4884 5101 5087 1 5079 2 AOI22S $T=929380 638520 1 180 $X=925660 $Y=638140
X2777 4963 5021 5119 5125 1 5132 2 AOI22S $T=926900 658680 0 0 $X=926900 $Y=658300
X2778 5007 5103 5161 5113 1 5134 2 AOI22S $T=934960 699000 1 180 $X=931240 $Y=698620
X2779 5153 991 5140 5107 1 5173 2 AOI22S $T=933720 588120 1 0 $X=933720 $Y=582700
X2780 5170 5021 5172 5163 1 5160 2 AOI22S $T=937440 658680 0 180 $X=933720 $Y=653260
X2781 5153 991 5165 5174 1 5179 2 AOI22S $T=934960 567960 1 0 $X=934960 $Y=562540
X2782 5153 991 5136 5148 1 993 2 AOI22S $T=935580 547800 1 0 $X=935580 $Y=542380
X2783 5170 991 5024 5178 1 5177 2 AOI22S $T=935580 598200 1 0 $X=935580 $Y=592780
X2784 5091 5159 5164 5157 1 5168 2 AOI22S $T=935580 638520 0 0 $X=935580 $Y=638140
X2785 5153 991 5150 5182 1 5192 2 AOI22S $T=936200 547800 0 0 $X=936200 $Y=547420
X2786 5102 5089 5166 5193 1 5184 2 AOI22S $T=937440 678840 1 0 $X=937440 $Y=673420
X2787 5170 5196 5158 5199 1 5128 2 AOI22S $T=938680 608280 1 0 $X=938680 $Y=602860
X2788 5102 5089 5211 5227 1 5237 2 AOI22S $T=943640 678840 1 0 $X=943640 $Y=673420
X2789 5007 5103 5222 5231 1 5202 2 AOI22S $T=943640 699000 1 0 $X=943640 $Y=693580
X2790 5007 5103 5212 5228 1 5238 2 AOI22S $T=943640 699000 0 0 $X=943640 $Y=698620
X2791 5102 5089 5226 5233 1 5232 2 AOI22S $T=944260 688920 1 0 $X=944260 $Y=683500
X2792 998 999 5121 1002 1 1001 2 AOI22S $T=945500 547800 1 0 $X=945500 $Y=542380
X2793 5214 1000 5123 5251 1 5249 2 AOI22S $T=951700 588120 0 180 $X=947980 $Y=582700
X2794 4963 5217 5247 5258 1 5254 2 AOI22S $T=948600 658680 0 0 $X=948600 $Y=658300
X2795 5214 999 5138 1003 1 1004 2 AOI22S $T=949220 547800 1 0 $X=949220 $Y=542380
X2796 4963 5217 5245 5269 1 5265 2 AOI22S $T=949840 668760 1 0 $X=949840 $Y=663340
X2797 5091 5261 5225 5253 1 1005 2 AOI22S $T=950460 638520 0 0 $X=950460 $Y=638140
X2798 5214 1000 5122 5282 1 5270 2 AOI22S $T=951700 567960 1 0 $X=951700 $Y=562540
X2799 5091 1000 5142 5289 1 1010 2 AOI22S $T=953560 618360 1 0 $X=953560 $Y=612940
X2800 5214 1000 5041 5293 1 5302 2 AOI22S $T=954800 608280 1 0 $X=954800 $Y=602860
X2801 5214 1000 5002 5316 1 5328 2 AOI22S $T=960380 608280 0 0 $X=960380 $Y=607900
X2802 5424 5403 5419 5391 1 5398 2 AOI22S $T=984560 699000 0 180 $X=980840 $Y=693580
X2803 5422 5402 5413 5409 1 5367 2 AOI22S $T=985800 658680 0 180 $X=982080 $Y=653260
X2804 5422 5402 5423 5397 1 5377 2 AOI22S $T=987040 668760 1 180 $X=983320 $Y=668380
X2805 5424 5403 5444 5404 1 5387 2 AOI22S $T=990760 578040 1 180 $X=987040 $Y=577660
X2806 1056 1051 5427 5338 1 5342 2 AOI22S $T=990760 598200 1 180 $X=987040 $Y=597820
X2807 1056 1051 5433 5380 1 5384 2 AOI22S $T=990760 628440 1 180 $X=987040 $Y=628060
X2808 5428 1052 5451 1050 1 1035 2 AOI22S $T=991380 547800 0 180 $X=987660 $Y=542380
X2809 5455 5460 5439 5431 1 5472 2 AOI22S $T=990140 668760 1 0 $X=990140 $Y=663340
X2810 1056 1051 5491 5476 1 5432 2 AOI22S $T=995720 598200 1 180 $X=992000 $Y=597820
X2811 5424 5403 5473 5462 1 5447 2 AOI22S $T=992620 688920 0 0 $X=992620 $Y=688540
X2812 5512 5446 5481 5487 1 5381 2 AOI22S $T=999440 638520 0 180 $X=995720 $Y=633100
X2813 5483 5496 5490 5500 1 5468 2 AOI22S $T=995720 658680 0 0 $X=995720 $Y=658300
X2814 5502 1052 5520 1065 1 5410 2 AOI22S $T=1000060 557880 0 180 $X=996340 $Y=552460
X2815 5483 5496 5426 5509 1 5515 2 AOI22S $T=997580 608280 1 0 $X=997580 $Y=602860
X2816 1056 1082 5523 5336 1 5514 2 AOI22S $T=1001300 547800 0 0 $X=1001300 $Y=547420
X2817 5455 5460 5526 5548 1 5550 2 AOI22S $T=1003780 668760 1 0 $X=1003780 $Y=663340
X2818 5512 5446 5527 5530 1 5540 2 AOI22S $T=1004400 638520 1 0 $X=1004400 $Y=633100
X2819 5545 5554 5544 5533 1 5562 2 AOI22S $T=1005020 699000 1 0 $X=1005020 $Y=693580
X2820 1087 1088 5506 5588 1 1089 2 AOI22S $T=1009980 547800 0 0 $X=1009980 $Y=547420
X2821 1087 1088 5573 5565 1 5583 2 AOI22S $T=1010600 557880 0 0 $X=1010600 $Y=557500
X2822 5568 1088 5435 5558 1 5599 2 AOI22S $T=1011220 578040 1 0 $X=1011220 $Y=572620
X2823 5422 5402 5537 5592 1 5600 2 AOI22S $T=1011220 588120 0 0 $X=1011220 $Y=587740
X2824 5422 5589 5538 5594 1 5572 2 AOI22S $T=1011220 668760 0 0 $X=1011220 $Y=668380
X2825 5455 5460 5627 5615 1 5634 2 AOI22S $T=1016180 658680 0 0 $X=1016180 $Y=658300
X2826 5545 5554 5633 5628 1 5602 2 AOI22S $T=1019900 699000 0 180 $X=1016180 $Y=693580
X2827 5512 5446 5632 5585 1 5655 2 AOI22S $T=1019900 638520 1 0 $X=1019900 $Y=633100
X2828 5672 5589 5642 5640 1 5641 2 AOI22S $T=1026100 668760 1 180 $X=1022380 $Y=668380
X2829 5543 1103 5561 5665 1 1105 2 AOI22S $T=1023000 557880 0 0 $X=1023000 $Y=557500
X2830 5543 1103 5497 5679 1 1106 2 AOI22S $T=1024860 537720 0 0 $X=1024860 $Y=537340
X2831 5681 5460 5687 5684 1 5678 2 AOI22S $T=1028580 658680 0 0 $X=1028580 $Y=658300
X2832 5512 5446 5715 5700 1 5698 2 AOI22S $T=1032920 618360 0 180 $X=1029200 $Y=612940
X2833 5512 5446 5692 5667 1 5636 2 AOI22S $T=1032920 628440 1 180 $X=1029200 $Y=628060
X2834 5545 5554 5704 5657 1 5688 2 AOI22S $T=1032920 688920 1 180 $X=1029200 $Y=688540
X2835 5672 5589 5701 5685 1 5719 2 AOI22S $T=1032920 668760 1 0 $X=1032920 $Y=663340
X2836 5545 5554 5735 5736 1 5742 2 AOI22S $T=1036640 688920 0 0 $X=1036640 $Y=688540
X2837 5762 5745 5716 5689 1 5738 2 AOI22S $T=1041600 608280 0 180 $X=1037880 $Y=602860
X2838 5720 5744 5725 5663 1 5669 2 AOI22S $T=1038500 578040 1 0 $X=1038500 $Y=572620
X2839 5672 5589 5746 5737 1 5753 2 AOI22S $T=1039120 668760 1 0 $X=1039120 $Y=663340
X2840 5762 5745 5775 5749 1 5764 2 AOI22S $T=1044700 598200 1 0 $X=1044700 $Y=592780
X2841 5720 5744 5792 5785 1 5743 2 AOI22S $T=1050280 578040 0 180 $X=1046560 $Y=572620
X2842 5518 5755 5827 5454 1 5811 2 AOI22S $T=1055240 628440 1 180 $X=1051520 $Y=628060
X2843 5502 5777 5810 5824 1 5814 2 AOI22S $T=1052140 557880 0 0 $X=1052140 $Y=557500
X2844 5693 5589 5825 5754 1 5837 2 AOI22S $T=1053380 668760 1 0 $X=1053380 $Y=663340
X2845 5829 5554 5849 5833 1 5839 2 AOI22S $T=1059580 688920 1 180 $X=1055860 $Y=688540
X2846 5868 5861 5801 5847 1 5856 2 AOI22S $T=1062680 598200 0 180 $X=1058960 $Y=592780
X2847 5681 5817 5840 5773 1 5823 2 AOI22S $T=1059580 668760 0 0 $X=1059580 $Y=668380
X2848 5502 5777 5874 5646 1 5846 2 AOI22S $T=1063300 557880 0 0 $X=1063300 $Y=557500
X2849 5868 5861 5859 5885 1 5843 2 AOI22S $T=1063920 588120 0 0 $X=1063920 $Y=587740
X2850 5868 5861 5904 5927 1 5867 2 AOI22S $T=1068260 588120 0 0 $X=1068260 $Y=587740
X2851 5681 5817 5891 5879 1 5929 2 AOI22S $T=1070740 678840 0 0 $X=1070740 $Y=678460
X2852 5720 5744 5933 5908 1 1147 2 AOI22S $T=1075080 567960 0 0 $X=1075080 $Y=567580
X2853 5935 5777 5940 1151 1 5961 2 AOI22S $T=1076940 547800 0 0 $X=1076940 $Y=547420
X2854 5681 5817 5973 5960 1 5938 2 AOI22S $T=1083140 678840 1 180 $X=1079420 $Y=678460
X2855 5680 5745 5921 5949 1 5968 2 AOI22S $T=1080040 598200 1 0 $X=1080040 $Y=592780
X2856 5981 5817 5982 5977 1 5939 2 AOI22S $T=1086860 658680 1 180 $X=1083140 $Y=658300
X2857 5680 5994 5999 5986 1 5990 2 AOI22S $T=1089340 588120 0 180 $X=1085620 $Y=582700
X2858 5981 5817 6015 5943 1 5969 2 AOI22S $T=1091200 658680 1 180 $X=1087480 $Y=658300
X2859 5981 5817 6029 6007 1 5988 2 AOI22S $T=1093680 668760 0 180 $X=1089960 $Y=663340
X2860 6008 5996 6024 6000 1 5953 2 AOI22S $T=1094300 628440 1 180 $X=1090580 $Y=628060
X2861 5829 5682 6038 6034 1 5978 2 AOI22S $T=1096780 699000 1 180 $X=1093060 $Y=698620
X2862 6008 5996 6012 6041 1 5979 2 AOI22S $T=1094300 628440 0 0 $X=1094300 $Y=628060
X2863 5935 6016 6053 1165 1 6022 2 AOI22S $T=1098640 557880 1 180 $X=1094920 $Y=557500
X2864 5680 5745 6055 6009 1 6037 2 AOI22S $T=1098640 608280 0 180 $X=1094920 $Y=602860
X2865 5829 5682 6058 6049 1 6003 2 AOI22S $T=1099260 699000 0 180 $X=1095540 $Y=693580
X2866 6008 5996 6045 6043 1 5974 2 AOI22S $T=1096160 638520 1 0 $X=1096160 $Y=633100
X2867 5935 6016 6062 1173 1 6070 2 AOI22S $T=1098640 557880 0 0 $X=1098640 $Y=557500
X2868 5829 5682 6051 6069 1 6071 2 AOI22S $T=1099260 699000 1 0 $X=1099260 $Y=693580
X2869 5518 5996 6068 6082 1 6073 2 AOI22S $T=1101120 638520 1 0 $X=1101120 $Y=633100
X2870 5693 5911 6074 6107 1 6108 2 AOI22S $T=1104220 618360 1 0 $X=1104220 $Y=612940
X2871 5720 6110 6023 6113 1 1180 2 AOI22S $T=1105460 557880 0 0 $X=1105460 $Y=557500
X2872 6104 5996 6100 6119 1 6103 2 AOI22S $T=1106080 608280 1 0 $X=1106080 $Y=602860
X2873 6118 5911 6042 6133 1 6129 2 AOI22S $T=1107940 668760 1 0 $X=1107940 $Y=663340
X2874 6118 5911 6079 6128 1 6139 2 AOI22S $T=1108560 658680 0 0 $X=1108560 $Y=658300
X2875 5720 6110 6067 6061 1 6142 2 AOI22S $T=1109180 557880 0 0 $X=1109180 $Y=557500
X2876 6104 5861 6064 6135 1 6160 2 AOI22S $T=1109180 588120 0 0 $X=1109180 $Y=587740
X2877 6118 5911 6057 6105 1 6143 2 AOI22S $T=1109180 668760 0 0 $X=1109180 $Y=668380
X2878 6118 5911 6019 6122 1 6149 2 AOI22S $T=1109800 678840 1 0 $X=1109800 $Y=673420
X2879 3734 3737 3688 3729 2 1 3764 AN4S $T=673320 668760 0 0 $X=673320 $Y=668380
X2880 3802 3782 3673 3813 2 1 3825 AN4S $T=685720 588120 0 0 $X=685720 $Y=587740
X2881 3808 3810 3618 3758 2 1 3828 AN4S $T=686960 658680 1 0 $X=686960 $Y=653260
X2882 3801 3812 3619 3795 2 1 3833 AN4S $T=687580 668760 1 0 $X=687580 $Y=663340
X2883 3789 3818 3617 3830 2 1 3865 AN4S $T=689440 567960 1 0 $X=689440 $Y=562540
X2884 3794 3784 3745 3835 2 1 3848 AN4S $T=690060 557880 1 0 $X=690060 $Y=552460
X2885 3852 3854 3651 3857 2 1 3874 AN4S $T=694400 678840 1 0 $X=694400 $Y=673420
X2886 3817 3895 3674 3899 2 1 3909 AN4S $T=702460 567960 1 0 $X=702460 $Y=562540
X2887 3908 3869 3675 3921 2 1 3931 AN4S $T=708660 598200 0 0 $X=708660 $Y=597820
X2888 3910 3915 3638 3919 2 1 3939 AN4S $T=709900 658680 0 0 $X=709900 $Y=658300
X2889 3977 3987 3991 3983 2 1 4009 AN4S $T=723540 608280 1 0 $X=723540 $Y=602860
X2890 3981 3994 3982 4004 2 1 4017 AN4S $T=724780 668760 0 0 $X=724780 $Y=668380
X2891 4152 4147 4146 4182 2 1 4190 AN4S $T=757640 608280 0 0 $X=757640 $Y=607900
X2892 4166 4202 4206 4211 2 1 4222 AN4S $T=763840 678840 0 0 $X=763840 $Y=678460
X2893 4088 4231 4215 4241 2 1 4248 AN4S $T=769420 598200 0 0 $X=769420 $Y=597820
X2894 4172 4267 4224 4276 2 1 4288 AN4S $T=776860 578040 1 0 $X=776860 $Y=572620
X2895 4186 4272 4263 4286 2 1 4307 AN4S $T=779340 658680 0 0 $X=779340 $Y=658300
X2896 4151 4297 4306 4311 2 1 4323 AN4S $T=783060 578040 1 0 $X=783060 $Y=572620
X2897 4161 4298 4303 4312 2 1 4324 AN4S $T=783060 588120 0 0 $X=783060 $Y=587740
X2898 4189 4309 4314 4322 2 1 4332 AN4S $T=784920 668760 0 0 $X=784920 $Y=668380
X2899 4098 4336 4346 4350 2 1 4359 AN4S $T=791120 678840 1 0 $X=791120 $Y=673420
X2900 4163 4364 4369 4368 2 1 4403 AN4S $T=798560 668760 0 0 $X=798560 $Y=668380
X2901 4154 4372 4302 4363 2 1 4421 AN4S $T=802280 567960 0 0 $X=802280 $Y=567580
X2902 4081 4392 4374 4391 2 1 4430 AN4S $T=804760 658680 0 0 $X=804760 $Y=658300
X2903 4533 4527 4516 4510 2 1 4474 AN4S $T=828320 668760 1 180 $X=823360 $Y=668380
X2904 4602 4593 4589 4586 2 1 4480 AN4S $T=838860 668760 0 180 $X=833900 $Y=663340
X2905 4616 4584 4618 4611 2 1 4507 AN4S $T=843820 588120 1 180 $X=838860 $Y=587740
X2906 4596 4648 4641 4640 2 1 4497 AN4S $T=847540 658680 0 180 $X=842580 $Y=653260
X2907 4646 4597 4647 4644 2 1 4470 AN4S $T=848780 557880 0 180 $X=843820 $Y=552460
X2908 4628 4600 4642 4649 2 1 4471 AN4S $T=843820 598200 0 0 $X=843820 $Y=597820
X2909 4667 4587 4680 4687 2 1 4447 AN4S $T=850640 567960 0 0 $X=850640 $Y=567580
X2910 4698 4700 4721 4729 2 1 4699 AN4S $T=856220 668760 0 0 $X=856220 $Y=668380
X2911 4629 4750 4771 4777 2 1 4758 AN4S $T=865520 668760 0 0 $X=865520 $Y=668380
X2912 4872 4861 4853 4843 2 1 4493 AN4S $T=884120 678840 0 180 $X=879160 $Y=673420
X2913 4991 4980 4972 4970 2 1 4454 AN4S $T=905200 678840 0 180 $X=900240 $Y=673420
X2914 4997 4988 4981 4965 2 1 4437 AN4S $T=906440 678840 1 180 $X=901480 $Y=678460
X2915 5024 4934 5005 5002 2 1 4531 AN4S $T=910160 608280 0 180 $X=905200 $Y=602860
X2916 5054 4975 5043 5041 2 1 4501 AN4S $T=915740 608280 1 180 $X=910780 $Y=607900
X2917 5119 5093 5106 5101 2 1 4434 AN4S $T=927520 678840 0 180 $X=922560 $Y=673420
X2918 5136 5019 5064 5121 2 1 5108 AN4S $T=930620 547800 0 180 $X=925660 $Y=542380
X2919 5150 4982 5074 5122 2 1 5105 AN4S $T=930620 557880 0 180 $X=925660 $Y=552460
X2920 5140 4992 5086 5123 2 1 5112 AN4S $T=930620 588120 0 180 $X=925660 $Y=582700
X2921 5165 4994 5083 5138 2 1 5030 AN4S $T=933720 567960 0 180 $X=928760 $Y=562540
X2922 5158 4908 5065 5142 2 1 5124 AN4S $T=934340 618360 0 180 $X=929380 $Y=612940
X2923 5172 5161 5166 5164 2 1 4460 AN4S $T=937440 658680 1 180 $X=932480 $Y=658300
X2924 5245 5222 5211 5225 2 1 4440 AN4S $T=947980 658680 1 180 $X=943020 $Y=658300
X2925 5247 5212 5226 5230 2 1 4452 AN4S $T=948600 668760 1 180 $X=943640 $Y=668380
X2926 5444 5435 5427 5426 2 1 5117 AN4S $T=988900 588120 1 180 $X=983940 $Y=587740
X2927 5419 5423 5433 5439 2 1 4490 AN4S $T=985180 668760 1 0 $X=985180 $Y=663340
X2928 5473 5413 5481 5490 2 1 4489 AN4S $T=992620 658680 1 0 $X=992620 $Y=653260
X2929 5451 5506 1077 5497 2 1 5023 AN4S $T=1000060 547800 0 180 $X=995100 $Y=542380
X2930 5511 5537 5491 5524 2 1 4526 AN4S $T=1005020 598200 1 180 $X=1000060 $Y=597820
X2931 5544 5538 5527 5526 2 1 4695 AN4S $T=1005020 668760 1 180 $X=1000060 $Y=668380
X2932 5520 5573 5523 5561 2 1 5097 AN4S $T=1010600 557880 1 180 $X=1005640 $Y=557500
X2933 5633 5642 5632 5627 2 1 4472 AN4S $T=1021140 668760 1 180 $X=1016180 $Y=668380
X2934 5704 5701 5692 5687 2 1 4748 AN4S $T=1031680 668760 1 180 $X=1026720 $Y=668380
X2935 5730 5725 5715 5716 2 1 4498 AN4S $T=1037260 608280 0 180 $X=1032300 $Y=602860
X2936 5735 5746 5741 5739 2 1 4475 AN4S $T=1041600 678840 0 180 $X=1036640 $Y=673420
X2937 5810 5792 5801 5775 2 1 5118 AN4S $T=1052760 588120 1 180 $X=1047800 $Y=587740
X2938 5874 5864 5859 5855 2 1 4504 AN4S $T=1062680 588120 1 180 $X=1057720 $Y=587740
X2939 5880 5899 5878 5891 2 1 4449 AN4S $T=1068880 678840 1 180 $X=1063920 $Y=678460
X2940 5940 5933 5904 5921 2 1 4445 AN4S $T=1075700 578040 0 180 $X=1070740 $Y=572620
X2941 6027 6019 6012 5973 2 1 4433 AN4S $T=1093680 678840 0 180 $X=1088720 $Y=673420
X2942 6030 6023 6014 5999 2 1 4466 AN4S $T=1094300 588120 0 180 $X=1089340 $Y=582700
X2943 6051 6042 6024 6015 2 1 4438 AN4S $T=1097400 658680 1 180 $X=1092440 $Y=658300
X2944 6038 6057 6045 6029 2 1 4451 AN4S $T=1099260 668760 0 180 $X=1094300 $Y=663340
X2945 6062 6067 6064 6044 2 1 4513 AN4S $T=1102360 578040 1 180 $X=1097400 $Y=577660
X2946 6058 6079 6068 5982 2 1 4455 AN4S $T=1103600 658680 1 180 $X=1098640 $Y=658300
X2947 6100 6055 6074 6053 2 1 4467 AN4S $T=1104220 608280 0 180 $X=1099260 $Y=602860
X2948 1491 2 1 54 BUF1 $T=265980 547800 0 180 $X=263500 $Y=542380
X2949 1543 2 1 1421 BUF1 $T=274040 668760 0 0 $X=274040 $Y=668380
X2950 1551 2 1 72 BUF1 $T=282100 537720 1 180 $X=279620 $Y=537340
X2951 1578 2 1 1551 BUF1 $T=282720 547800 0 0 $X=282720 $Y=547420
X2952 1656 2 1 1455 BUF1 $T=301320 668760 1 180 $X=298840 $Y=668380
X2953 1641 2 1 1675 BUF1 $T=303180 567960 0 0 $X=303180 $Y=567580
X2954 1703 2 1 79 BUF1 $T=306280 678840 1 180 $X=303800 $Y=678460
X2955 1816 2 1 1770 BUF1 $T=325500 557880 1 0 $X=325500 $Y=552460
X2956 1701 2 1 1835 BUF1 $T=325500 668760 1 0 $X=325500 $Y=663340
X2957 148 2 1 121 BUF1 $T=337280 567960 1 180 $X=334800 $Y=567580
X2958 1876 2 1 1733 BUF1 $T=340380 547800 1 180 $X=337900 $Y=547420
X2959 1858 2 1 1905 BUF1 $T=342860 578040 0 0 $X=342860 $Y=577660
X2960 1864 2 1 1930 BUF1 $T=349680 678840 0 0 $X=349680 $Y=678460
X2961 1864 2 1 1982 BUF1 $T=362080 608280 0 0 $X=362080 $Y=607900
X2962 1612 2 1 2039 BUF1 $T=369520 567960 0 0 $X=369520 $Y=567580
X2963 2066 2 1 2065 BUF1 $T=373240 567960 0 0 $X=373240 $Y=567580
X2964 2239 2 1 210 BUF1 $T=411060 588120 0 180 $X=408580 $Y=582700
X2965 2277 2 1 234 BUF1 $T=419740 719160 0 0 $X=419740 $Y=718780
X2966 2357 2 1 211 BUF1 $T=425940 588120 0 180 $X=423460 $Y=582700
X2967 148 2 1 2410 BUF1 $T=437100 578040 0 0 $X=437100 $Y=577660
X2968 2504 2 1 2387 BUF1 $T=452600 638520 1 180 $X=450120 $Y=638140
X2969 2583 2 1 271 BUF1 $T=465000 598200 0 180 $X=462520 $Y=592780
X2970 2658 2 1 275 BUF1 $T=478640 547800 1 180 $X=476160 $Y=547420
X2971 2687 2 1 2668 BUF1 $T=487940 588120 1 180 $X=485460 $Y=587740
X2972 331 2 1 2687 BUF1 $T=501580 588120 1 180 $X=499100 $Y=587740
X2973 2790 2 1 2741 BUF1 $T=500340 638520 0 0 $X=500340 $Y=638140
X2974 295 2 1 2729 BUF1 $T=507160 588120 1 180 $X=504680 $Y=587740
X2975 2889 2 1 2868 BUF1 $T=521420 709080 1 180 $X=518940 $Y=708700
X2976 2962 2 1 2858 BUF1 $T=530100 719160 0 180 $X=527620 $Y=713740
X2977 346 2 1 2614 BUF1 $T=541260 578040 1 0 $X=541260 $Y=572620
X2978 433 2 1 2889 BUF1 $T=560480 709080 1 180 $X=558000 $Y=708700
X2979 425 2 1 3203 BUF1 $T=571640 547800 1 0 $X=571640 $Y=542380
X2980 473 2 1 413 BUF1 $T=576600 547800 0 180 $X=574120 $Y=542380
X2981 3192 2 1 2633 BUF1 $T=580320 588120 0 180 $X=577840 $Y=582700
X2982 437 2 1 3218 BUF1 $T=581560 588120 1 0 $X=581560 $Y=582700
X2983 343 2 1 3284 BUF1 $T=590240 709080 0 0 $X=590240 $Y=708700
X2984 3155 2 1 537 BUF1 $T=601400 578040 1 0 $X=601400 $Y=572620
X2985 473 2 1 3350 BUF1 $T=606360 537720 0 0 $X=606360 $Y=537340
X2986 406 2 1 3364 BUF1 $T=606980 578040 1 0 $X=606980 $Y=572620
X2987 512 2 1 3363 BUF1 $T=609460 547800 0 0 $X=609460 $Y=547420
X2988 3070 2 1 552 BUF1 $T=613180 567960 0 180 $X=610700 $Y=562540
X2989 40 2 1 3414 BUF1 $T=616280 699000 0 0 $X=616280 $Y=698620
X2990 542 2 1 3423 BUF1 $T=616900 688920 1 0 $X=616900 $Y=683500
X2991 3159 2 1 3613 BUF1 $T=650380 688920 0 0 $X=650380 $Y=688540
X2992 3544 2 1 3603 BUF1 $T=655960 628440 0 0 $X=655960 $Y=628060
X2993 3654 2 1 3607 BUF1 $T=660920 618360 0 180 $X=658440 $Y=612940
X2994 3660 2 1 3615 BUF1 $T=663400 668760 1 180 $X=660920 $Y=668380
X2995 3544 2 1 656 BUF1 $T=662160 699000 0 0 $X=662160 $Y=698620
X2996 3613 2 1 3665 BUF1 $T=662780 658680 0 0 $X=662780 $Y=658300
X2997 3654 2 1 661 BUF1 $T=664640 588120 1 0 $X=664640 $Y=582700
X2998 3665 2 1 3708 BUF1 $T=666500 588120 0 0 $X=666500 $Y=587740
X2999 3728 2 1 3654 BUF1 $T=672700 608280 0 180 $X=670220 $Y=602860
X3000 3708 2 1 669 BUF1 $T=672700 557880 1 0 $X=672700 $Y=552460
X3001 3537 2 1 3738 BUF1 $T=673320 628440 0 0 $X=673320 $Y=628060
X3002 3786 2 1 680 BUF1 $T=684480 567960 1 0 $X=684480 $Y=562540
X3003 3820 2 1 681 BUF1 $T=688820 578040 1 180 $X=686340 $Y=577660
X3004 3458 2 1 3832 BUF1 $T=691300 678840 1 0 $X=691300 $Y=673420
X3005 701 2 1 704 BUF1 $T=698740 537720 0 0 $X=698740 $Y=537340
X3006 3738 2 1 698 BUF1 $T=701220 567960 0 180 $X=698740 $Y=562540
X3007 705 2 1 3788 BUF1 $T=704320 598200 1 180 $X=701840 $Y=597820
X3008 703 2 1 3658 BUF1 $T=701840 668760 1 0 $X=701840 $Y=663340
X3009 3692 2 1 3902 BUF1 $T=703080 688920 1 0 $X=703080 $Y=683500
X3010 3658 2 1 701 BUF1 $T=708660 618360 1 0 $X=708660 $Y=612940
X3011 3951 2 1 715 BUF1 $T=716100 598200 0 0 $X=716100 $Y=597820
X3012 3562 2 1 3958 BUF1 $T=716100 668760 0 0 $X=716100 $Y=668380
X3013 3958 2 1 3951 BUF1 $T=717340 638520 0 0 $X=717340 $Y=638140
X3014 3888 2 1 721 BUF1 $T=717960 557880 0 0 $X=717960 $Y=557500
X3015 3996 2 1 3786 BUF1 $T=726640 598200 0 180 $X=724160 $Y=592780
X3016 4019 2 1 732 BUF1 $T=729740 557880 1 0 $X=729740 $Y=552460
X3017 4019 2 1 3820 BUF1 $T=732220 588120 0 0 $X=732220 $Y=587740
X3018 716 2 1 4068 BUF1 $T=740280 658680 0 0 $X=740280 $Y=658300
X3019 4080 2 1 4019 BUF1 $T=743380 648600 0 180 $X=740900 $Y=643180
X3020 4111 2 1 4116 BUF1 $T=747100 648600 1 0 $X=747100 $Y=643180
X3021 770 2 1 772 BUF1 $T=750200 699000 1 0 $X=750200 $Y=693580
X3022 3978 2 1 3996 BUF1 $T=758260 658680 0 0 $X=758260 $Y=658300
X3023 763 2 1 4157 BUF1 $T=758880 668760 1 0 $X=758880 $Y=663340
X3024 4180 2 1 3979 BUF1 $T=761360 678840 0 180 $X=758880 $Y=673420
X3025 4176 2 1 3992 BUF1 $T=759500 618360 1 0 $X=759500 $Y=612940
X3026 663 2 1 4173 BUF1 $T=762600 638520 1 0 $X=762600 $Y=633100
X3027 4173 2 1 748 BUF1 $T=764460 598200 1 0 $X=764460 $Y=592780
X3028 790 2 1 4184 BUF1 $T=766940 709080 1 180 $X=764460 $Y=708700
X3029 457 2 1 4223 BUF1 $T=764460 719160 0 0 $X=764460 $Y=718780
X3030 3979 2 1 793 BUF1 $T=767560 578040 1 0 $X=767560 $Y=572620
X3031 3979 2 1 3728 BUF1 $T=770660 608280 1 180 $X=768180 $Y=607900
X3032 3660 2 1 4218 BUF1 $T=769420 678840 0 0 $X=769420 $Y=678460
X3033 4168 2 1 4254 BUF1 $T=773140 628440 0 0 $X=773140 $Y=628060
X3034 4148 2 1 4258 BUF1 $T=773760 638520 1 0 $X=773760 $Y=633100
X3035 678 2 1 4253 BUF1 $T=782440 668760 0 0 $X=782440 $Y=668380
X3036 3992 2 1 808 BUF1 $T=784300 578040 0 0 $X=784300 $Y=577660
X3037 802 2 1 4188 BUF1 $T=787400 537720 1 180 $X=784920 $Y=537340
X3038 3701 2 1 816 BUF1 $T=788020 638520 1 0 $X=788020 $Y=633100
X3039 4343 2 1 802 BUF1 $T=791120 537720 1 180 $X=788640 $Y=537340
X3040 4067 2 1 4233 BUF1 $T=789880 668760 0 0 $X=789880 $Y=668380
X3041 4233 2 1 814 BUF1 $T=792980 578040 1 0 $X=792980 $Y=572620
X3042 4025 2 1 801 BUF1 $T=793600 598200 0 0 $X=793600 $Y=597820
X3043 4106 2 1 798 BUF1 $T=794840 537720 0 0 $X=794840 $Y=537340
X3044 818 2 1 822 BUF1 $T=797940 557880 0 0 $X=797940 $Y=557500
X3045 4068 2 1 4343 BUF1 $T=804760 618360 0 0 $X=804760 $Y=617980
X3046 4068 2 1 4423 BUF1 $T=806000 678840 1 0 $X=806000 $Y=673420
X3047 4183 2 1 4537 BUF1 $T=821500 598200 0 0 $X=821500 $Y=597820
X3048 4253 2 1 4515 BUF1 $T=822740 628440 1 0 $X=822740 $Y=623020
X3049 4343 2 1 863 BUF1 $T=827080 567960 0 0 $X=827080 $Y=567580
X3050 849 2 1 4582 BUF1 $T=834520 638520 1 0 $X=834520 $Y=633100
X3051 4583 2 1 4591 BUF1 $T=835140 658680 1 0 $X=835140 $Y=653260
X3052 4588 2 1 4573 BUF1 $T=837000 638520 0 0 $X=837000 $Y=638140
X3053 4588 2 1 885 BUF1 $T=847540 567960 0 0 $X=847540 $Y=567580
X3054 4537 2 1 4674 BUF1 $T=849400 598200 0 0 $X=849400 $Y=597820
X3055 4534 2 1 4679 BUF1 $T=850020 699000 1 0 $X=850020 $Y=693580
X3056 4523 2 1 4692 BUF1 $T=851260 699000 0 0 $X=851260 $Y=698620
X3057 4591 2 1 895 BUF1 $T=853740 578040 1 0 $X=853740 $Y=572620
X3058 4561 2 1 4703 BUF1 $T=853740 668760 0 0 $X=853740 $Y=668380
X3059 863 2 1 4720 BUF1 $T=856840 567960 0 0 $X=856840 $Y=567580
X3060 4561 2 1 4718 BUF1 $T=856840 628440 1 0 $X=856840 $Y=623020
X3061 4719 2 1 4714 BUF1 $T=857460 648600 1 0 $X=857460 $Y=643180
X3062 819 2 1 4759 BUF1 $T=862420 709080 0 0 $X=862420 $Y=708700
X3063 892 2 1 4708 BUF1 $T=866140 588120 0 180 $X=863660 $Y=582700
X3064 4718 2 1 4786 BUF1 $T=866760 598200 1 0 $X=866760 $Y=592780
X3065 4477 2 1 917 BUF1 $T=868620 598200 0 0 $X=868620 $Y=597820
X3066 4500 2 1 919 BUF1 $T=869240 557880 0 0 $X=869240 $Y=557500
X3067 4477 2 1 4795 BUF1 $T=869860 648600 0 0 $X=869860 $Y=648220
X3068 4500 2 1 4803 BUF1 $T=874200 648600 1 0 $X=874200 $Y=643180
X3069 3902 2 1 4878 BUF1 $T=883500 628440 1 0 $X=883500 $Y=623020
X3070 4803 2 1 4884 BUF1 $T=883500 638520 0 0 $X=883500 $Y=638140
X3071 930 2 1 4900 BUF1 $T=886600 709080 0 0 $X=886600 $Y=708700
X3072 796 2 1 936 BUF1 $T=887840 719160 0 0 $X=887840 $Y=718780
X3073 873 2 1 4915 BUF1 $T=888460 567960 0 0 $X=888460 $Y=567580
X3074 4903 2 1 925 BUF1 $T=890940 598200 0 180 $X=888460 $Y=592780
X3075 4708 2 1 4912 BUF1 $T=889080 588120 1 0 $X=889080 $Y=582700
X3076 4583 2 1 4963 BUF1 $T=899620 658680 1 0 $X=899620 $Y=653260
X3077 4679 2 1 5007 BUF1 $T=903960 699000 1 0 $X=903960 $Y=693580
X3078 4714 2 1 947 BUF1 $T=905200 557880 1 0 $X=905200 $Y=552460
X3079 4573 2 1 5021 BUF1 $T=906440 658680 1 0 $X=906440 $Y=653260
X3080 4795 2 1 5091 BUF1 $T=918840 638520 0 0 $X=918840 $Y=638140
X3081 4714 2 1 974 BUF1 $T=919460 557880 1 0 $X=919460 $Y=552460
X3082 936 2 1 975 BUF1 $T=920080 719160 0 0 $X=920080 $Y=718780
X3083 4703 2 1 5089 BUF1 $T=920700 678840 0 0 $X=920700 $Y=678460
X3084 4692 2 1 5103 BUF1 $T=922560 699000 0 0 $X=922560 $Y=698620
X3085 938 2 1 968 BUF1 $T=922560 719160 0 0 $X=922560 $Y=718780
X3086 4515 2 1 965 BUF1 $T=926280 598200 1 180 $X=923800 $Y=597820
X3087 4903 2 1 985 BUF1 $T=927520 598200 1 0 $X=927520 $Y=592780
X3088 4515 2 1 5155 BUF1 $T=931240 608280 1 0 $X=931240 $Y=602860
X3089 4963 2 1 990 BUF1 $T=936200 628440 0 180 $X=933720 $Y=623020
X3090 4900 2 1 4903 BUF1 $T=940540 699000 0 0 $X=940540 $Y=698620
X3091 871 2 1 996 BUF1 $T=940540 719160 0 0 $X=940540 $Y=718780
X3092 5214 2 1 998 BUF1 $T=943020 547800 1 0 $X=943020 $Y=542380
X3093 974 2 1 5167 BUF1 $T=949220 557880 1 0 $X=949220 $Y=552460
X3094 4759 2 1 1017 BUF1 $T=957900 719160 0 0 $X=957900 $Y=718780
X3095 4423 2 1 5285 BUF1 $T=961620 678840 1 0 $X=961620 $Y=673420
X3096 5358 2 1 5100 BUF1 $T=973400 588120 1 0 $X=973400 $Y=582700
X3097 816 2 1 1034 BUF1 $T=978980 628440 1 0 $X=978980 $Y=623020
X3098 900 2 1 1046 BUF1 $T=984560 719160 1 0 $X=984560 $Y=713740
X3099 4969 2 1 5445 BUF1 $T=988280 608280 0 0 $X=988280 $Y=607900
X3100 4903 2 1 1058 BUF1 $T=988280 719160 1 0 $X=988280 $Y=713740
X3101 4630 2 1 1056 BUF1 $T=993860 638520 0 180 $X=991380 $Y=633100
X3102 5424 2 1 5502 BUF1 $T=993860 557880 1 0 $X=993860 $Y=552460
X3103 5482 2 1 5460 BUF1 $T=993860 668760 1 0 $X=993860 $Y=663340
X3104 5482 2 1 5496 BUF1 $T=996340 668760 1 0 $X=996340 $Y=663340
X3105 4630 2 1 5518 BUF1 $T=998200 628440 0 0 $X=998200 $Y=628060
X3106 5534 2 1 5424 BUF1 $T=1001300 688920 1 180 $X=998820 $Y=688540
X3107 5483 2 1 5543 BUF1 $T=1002540 608280 1 0 $X=1002540 $Y=602860
X3108 5483 2 1 5455 BUF1 $T=1002540 658680 0 0 $X=1002540 $Y=658300
X3109 5534 2 1 5545 BUF1 $T=1002540 688920 0 0 $X=1002540 $Y=688540
X3110 5402 2 1 1088 BUF1 $T=1008120 567960 0 0 $X=1008120 $Y=567580
X3111 1081 2 1 5519 BUF1 $T=1009360 699000 1 0 $X=1009360 $Y=693580
X3112 5402 2 1 5589 BUF1 $T=1011220 668760 1 0 $X=1011220 $Y=663340
X3113 5155 2 1 1097 BUF1 $T=1018040 608280 1 0 $X=1018040 $Y=602860
X3114 1097 2 1 5650 BUF1 $T=1019900 598200 0 0 $X=1019900 $Y=597820
X3115 5445 2 1 1101 BUF1 $T=1021760 588120 0 0 $X=1021760 $Y=587740
X3116 1086 2 1 5623 BUF1 $T=1023000 678840 0 0 $X=1023000 $Y=678460
X3117 5543 2 1 5680 BUF1 $T=1024240 588120 0 0 $X=1024240 $Y=587740
X3118 5496 2 1 1103 BUF1 $T=1026720 557880 0 0 $X=1026720 $Y=557500
X3119 5403 2 1 5682 BUF1 $T=1026720 688920 0 0 $X=1026720 $Y=688540
X3120 5422 2 1 5693 BUF1 $T=1027340 618360 0 0 $X=1027340 $Y=617980
X3121 1111 2 1 5674 BUF1 $T=1029200 678840 0 0 $X=1029200 $Y=678460
X3122 1090 2 1 5705 BUF1 $T=1032920 557880 0 0 $X=1032920 $Y=557500
X3123 5496 2 1 5745 BUF1 $T=1037880 598200 1 0 $X=1037880 $Y=592780
X3124 5680 2 1 5762 BUF1 $T=1041600 598200 1 0 $X=1041600 $Y=592780
X3125 1120 2 1 5777 BUF1 $T=1044700 557880 1 0 $X=1044700 $Y=552460
X3126 5446 2 1 5755 BUF1 $T=1044700 628440 0 0 $X=1044700 $Y=628060
X3127 1118 2 1 5781 BUF1 $T=1045940 709080 0 0 $X=1045940 $Y=708700
X3128 5797 2 1 1123 BUF1 $T=1050280 608280 0 0 $X=1050280 $Y=607900
X3129 5460 2 1 5817 BUF1 $T=1050900 668760 1 0 $X=1050900 $Y=663340
X3130 5545 2 1 5829 BUF1 $T=1052140 699000 1 0 $X=1052140 $Y=693580
X3131 5781 2 1 5797 BUF1 $T=1054620 678840 0 0 $X=1054620 $Y=678460
X3132 938 2 1 5858 BUF1 $T=1058960 719160 0 0 $X=1058960 $Y=718780
X3133 5518 2 1 5868 BUF1 $T=1060820 628440 0 0 $X=1060820 $Y=628060
X3134 938 2 1 1135 BUF1 $T=1063300 719160 0 0 $X=1063300 $Y=718780
X3135 4949 2 1 5897 BUF1 $T=1065160 638520 0 0 $X=1065160 $Y=638140
X3136 5589 2 1 5911 BUF1 $T=1068260 678840 1 0 $X=1068260 $Y=673420
X3137 1139 2 1 1142 BUF1 $T=1070120 719160 0 0 $X=1070120 $Y=718780
X3138 4949 2 1 1127 BUF1 $T=1071360 618360 1 0 $X=1071360 $Y=612940
X3139 5897 2 1 5890 BUF1 $T=1071360 668760 1 0 $X=1071360 $Y=663340
X3140 5502 2 1 5935 BUF1 $T=1072600 557880 0 0 $X=1072600 $Y=557500
X3141 1140 2 1 5946 BUF1 $T=1077560 598200 1 0 $X=1077560 $Y=592780
X3142 5890 2 1 1155 BUF1 $T=1081900 709080 1 0 $X=1081900 $Y=703660
X3143 5681 2 1 5981 BUF1 $T=1083140 668760 1 0 $X=1083140 $Y=663340
X3144 5755 2 1 5996 BUF1 $T=1085620 628440 0 0 $X=1085620 $Y=628060
X3145 5518 2 1 6008 BUF1 $T=1087480 628440 1 0 $X=1087480 $Y=623020
X3146 5732 2 1 5995 BUF1 $T=1088100 618360 1 0 $X=1088100 $Y=612940
X3147 5650 2 1 6013 BUF1 $T=1089340 638520 1 0 $X=1089340 $Y=633100
X3148 5745 2 1 5994 BUF1 $T=1093680 588120 0 0 $X=1093680 $Y=587740
X3149 5995 2 1 1164 BUF1 $T=1096780 557880 1 0 $X=1096780 $Y=552460
X3150 6005 2 1 6101 BUF1 $T=1104220 588120 0 0 $X=1104220 $Y=587740
X3151 5693 2 1 6118 BUF1 $T=1106080 668760 0 0 $X=1106080 $Y=668380
X3152 5996 2 1 5861 BUF1 $T=1106700 588120 0 0 $X=1106700 $Y=587740
X3153 5868 2 1 6104 BUF1 $T=1109800 598200 1 180 $X=1107320 $Y=597820
X3154 1156 2 1 6140 BUF1 $T=1109180 678840 0 0 $X=1109180 $Y=678460
X3155 6075 2 1 6056 BUF1 $T=1114140 618360 1 180 $X=1111660 $Y=617980
X3156 6140 2 1 6075 BUF1 $T=1116620 618360 1 180 $X=1114140 $Y=617980
X3157 1184 2 1 1146 BUF1 $T=1114140 719160 1 0 $X=1114140 $Y=713740
X3158 1270 1 2 1260 BUF1CK $T=223820 638520 1 0 $X=223820 $Y=633100
X3159 1275 1 2 1271 BUF1CK $T=224440 658680 1 0 $X=224440 $Y=653260
X3160 1280 1 2 1275 BUF1CK $T=225680 658680 0 0 $X=225680 $Y=658300
X3161 1284 1 2 1277 BUF1CK $T=226920 709080 0 0 $X=226920 $Y=708700
X3162 1287 1 2 1281 BUF1CK $T=230020 678840 0 0 $X=230020 $Y=678460
X3163 1369 1 2 1380 BUF1CK $T=244280 547800 1 0 $X=244280 $Y=542380
X3164 1576 1 2 1589 BUF1CK $T=281480 618360 0 0 $X=281480 $Y=617980
X3165 1703 1 2 1702 BUF1CK $T=306900 668760 0 180 $X=304420 $Y=663340
X3166 1656 1 2 1883 BUF1CK $T=342860 668760 1 0 $X=342860 $Y=663340
X3167 1896 1 2 1963 BUF1CK $T=352780 678840 1 0 $X=352780 $Y=673420
X3168 3597 1 2 3605 BUF1CK $T=652860 688920 0 0 $X=652860 $Y=688540
X3169 3528 1 2 3601 BUF1CK $T=655960 578040 0 0 $X=655960 $Y=577660
X3170 3709 1 2 3715 BUF1CK $T=667120 598200 0 0 $X=667120 $Y=597820
X3171 663 1 2 4169 BUF1CK $T=755780 709080 1 0 $X=755780 $Y=703660
X3172 4378 1 2 4387 BUF1CK $T=797940 699000 0 0 $X=797940 $Y=698620
X3173 4442 1 2 4450 BUF1CK $T=811580 719160 1 0 $X=811580 $Y=713740
X3174 830 1 2 832 BUF1CK $T=811580 719160 0 0 $X=811580 $Y=718780
X3175 4542 1 2 4517 BUF1CK $T=837620 688920 1 0 $X=837620 $Y=683500
X3176 4627 1 2 4632 BUF1CK $T=841960 719160 1 0 $X=841960 $Y=713740
X3177 4633 1 2 4639 BUF1CK $T=842580 638520 1 0 $X=842580 $Y=633100
X3178 4668 1 2 4671 BUF1CK $T=849400 608280 0 0 $X=849400 $Y=607900
X3179 4710 1 2 4722 BUF1CK $T=855600 709080 1 0 $X=855600 $Y=703660
X3180 4772 1 2 4779 BUF1CK $T=866760 648600 1 0 $X=866760 $Y=643180
X3181 4783 1 2 4768 BUF1CK $T=868620 678840 0 0 $X=868620 $Y=678460
X3182 4713 1 2 4737 BUF1CK $T=869240 638520 0 0 $X=869240 $Y=638140
X3183 4816 1 2 4766 BUF1CK $T=874820 688920 1 0 $X=874820 $Y=683500
X3184 4827 1 2 4849 BUF1CK $T=881020 588120 0 0 $X=881020 $Y=587740
X3185 4871 1 2 4869 BUF1CK $T=883500 668760 1 0 $X=883500 $Y=663340
X3186 4886 1 2 4895 BUF1CK $T=885980 678840 1 0 $X=885980 $Y=673420
X3187 4910 1 2 4815 BUF1CK $T=890940 628440 1 0 $X=890940 $Y=623020
X3188 4928 1 2 4933 BUF1CK $T=893420 557880 1 0 $X=893420 $Y=552460
X3189 4896 1 2 4890 BUF1CK $T=894660 699000 0 0 $X=894660 $Y=698620
X3190 4855 1 2 4836 BUF1CK $T=896520 608280 0 0 $X=896520 $Y=607900
X3191 4897 1 2 4825 BUF1CK $T=898380 638520 0 0 $X=898380 $Y=638140
X3192 4977 1 2 4983 BUF1CK $T=902720 578040 0 0 $X=902720 $Y=577660
X3193 4958 1 2 4961 BUF1CK $T=905200 688920 0 0 $X=905200 $Y=688540
X3194 5016 1 2 5025 BUF1CK $T=907680 648600 0 0 $X=907680 $Y=648220
X3195 5020 1 2 5009 BUF1CK $T=910160 608280 1 0 $X=910160 $Y=602860
X3196 5055 1 2 5016 BUF1CK $T=914500 648600 0 0 $X=914500 $Y=648220
X3197 5090 1 2 5057 BUF1CK $T=923180 557880 0 0 $X=923180 $Y=557500
X3198 5186 1 2 5195 BUF1CK $T=939920 547800 0 0 $X=939920 $Y=547420
X3199 5191 1 2 5218 BUF1CK $T=948600 668760 0 0 $X=948600 $Y=668380
X3200 5260 1 2 5246 BUF1CK $T=949840 588120 0 0 $X=949840 $Y=587740
X3201 5219 1 2 5274 BUF1CK $T=949840 709080 1 0 $X=949840 $Y=703660
X3202 5264 1 2 5236 BUF1CK $T=954800 598200 0 0 $X=954800 $Y=597820
X3203 1012 1 2 1014 BUF1CK $T=956040 709080 0 0 $X=956040 $Y=708700
X3204 5313 1 2 5310 BUF1CK $T=961000 658680 1 0 $X=961000 $Y=653260
X3205 5275 1 2 5235 BUF1CK $T=964720 598200 1 0 $X=964720 $Y=592780
X3206 5311 1 2 5319 BUF1CK $T=965340 567960 0 0 $X=965340 $Y=567580
X3207 5346 1 2 5357 BUF1CK $T=970920 699000 0 0 $X=970920 $Y=698620
X3208 5348 1 2 5356 BUF1CK $T=971540 688920 0 0 $X=971540 $Y=688540
X3209 5371 1 2 5376 BUF1CK $T=976500 658680 0 0 $X=976500 $Y=658300
X3210 5383 1 2 5392 BUF1CK $T=978980 547800 1 0 $X=978980 $Y=542380
X3211 5450 1 2 5459 BUF1CK $T=988900 678840 0 0 $X=988900 $Y=678460
X3212 5396 1 2 5429 BUF1CK $T=993860 628440 0 0 $X=993860 $Y=628060
X3213 1074 1 2 1069 BUF1CK $T=995100 537720 0 0 $X=995100 $Y=537340
X3214 5478 1 2 5486 BUF1CK $T=995100 598200 1 0 $X=995100 $Y=592780
X3215 5492 1 2 5479 BUF1CK $T=995720 719160 1 0 $X=995720 $Y=713740
X3216 5400 1 2 5437 BUF1CK $T=1000060 578040 0 0 $X=1000060 $Y=577660
X3217 5525 1 2 5529 BUF1CK $T=1001300 628440 0 0 $X=1001300 $Y=628060
X3218 5648 1 2 5635 BUF1CK $T=1020520 709080 1 0 $X=1020520 $Y=703660
X3219 1100 1 2 5586 BUF1CK $T=1022380 719160 0 0 $X=1022380 $Y=718780
X3220 5686 1 2 5677 BUF1CK $T=1029200 719160 1 0 $X=1029200 $Y=713740
X3221 5649 1 2 5631 BUF1CK $T=1032920 699000 1 0 $X=1032920 $Y=693580
X3222 5724 1 2 5733 BUF1CK $T=1034780 709080 1 0 $X=1034780 $Y=703660
X3223 5607 1 2 5690 BUF1CK $T=1035400 578040 0 0 $X=1035400 $Y=577660
X3224 5403 1 2 1120 BUF1CK $T=1039740 578040 0 0 $X=1039740 $Y=577660
X3225 5598 1 2 5604 BUF1CK $T=1040360 547800 0 0 $X=1040360 $Y=547420
X3226 5750 1 2 5761 BUF1CK $T=1040980 699000 0 0 $X=1040980 $Y=698620
X3227 5577 1 2 5643 BUF1CK $T=1042220 557880 1 0 $X=1042220 $Y=552460
X3228 1123 1 2 5760 BUF1CK $T=1044700 567960 1 0 $X=1044700 $Y=562540
X3229 5770 1 2 5800 BUF1CK $T=1049660 699000 1 0 $X=1049660 $Y=693580
X3230 5818 1 2 5828 BUF1CK $T=1052140 699000 0 0 $X=1052140 $Y=698620
X3231 5869 1 2 5876 BUF1CK $T=1061440 648600 0 0 $X=1061440 $Y=648220
X3232 5906 1 2 5901 BUF1CK $T=1068260 668760 0 0 $X=1068260 $Y=668380
X3233 5914 1 2 5913 BUF1CK $T=1070120 628440 1 0 $X=1070120 $Y=623020
X3234 5991 1 2 6010 BUF1CK $T=1088100 628440 0 0 $X=1088100 $Y=628060
X3235 5777 1 2 6016 BUF1CK $T=1089960 557880 1 0 $X=1089960 $Y=552460
X3236 5951 1 2 5930 BUF1CK $T=1091820 709080 1 0 $X=1091820 $Y=703660
X3237 6054 1 2 6060 BUF1CK $T=1097400 578040 1 0 $X=1097400 $Y=572620
X3238 6089 1 2 6096 BUF1CK $T=1102980 658680 1 0 $X=1102980 $Y=653260
X3239 6094 1 2 6151 BUF1CK $T=1125300 688920 0 0 $X=1125300 $Y=688540
X3240 6164 1 2 6112 BUF1CK $T=1126540 668760 1 0 $X=1126540 $Y=663340
X3241 1740 1703 1 2 INV2 $T=316820 678840 1 180 $X=314960 $Y=678460
X3242 1844 1701 1 2 INV2 $T=332320 648600 1 180 $X=330460 $Y=648220
X3243 2646 297 1 2 INV2 $T=476160 557880 0 0 $X=476160 $Y=557500
X3244 315 2630 1 2 INV2 $T=487940 557880 1 0 $X=487940 $Y=552460
X3245 346 2658 1 2 INV2 $T=507780 557880 0 0 $X=507780 $Y=557500
X3246 295 425 1 2 INV2 $T=554900 537720 0 0 $X=554900 $Y=537340
X3247 377 3155 1 2 INV2 $T=569160 537720 1 180 $X=567300 $Y=537340
X3248 415 3148 1 2 INV2 $T=567300 567960 0 0 $X=567300 $Y=567580
X3249 447 458 1 2 INV2 $T=569780 547800 1 0 $X=569780 $Y=542380
X3250 380 3182 1 2 INV2 $T=571020 567960 1 0 $X=571020 $Y=562540
X3251 378 474 1 2 INV2 $T=574740 557880 0 0 $X=574740 $Y=557500
X3252 437 3220 1 2 INV2 $T=597060 578040 1 0 $X=597060 $Y=572620
X3253 3687 3681 1 2 INV2 $T=664640 598200 0 0 $X=664640 $Y=597820
X3254 3873 3877 1 2 INV2 $T=698740 588120 0 0 $X=698740 $Y=587740
X3255 3892 702 1 2 INV2 $T=702460 557880 1 0 $X=702460 $Y=552460
X3256 4013 705 1 2 INV2 $T=728500 628440 0 0 $X=728500 $Y=628060
X3257 4013 4025 1 2 INV2 $T=730360 628440 0 0 $X=730360 $Y=628060
X3258 4062 708 1 2 INV2 $T=739660 618360 0 0 $X=739660 $Y=617980
X3259 4167 780 1 2 INV2 $T=759500 719160 1 0 $X=759500 $Y=713740
X3260 4594 4577 1 2 INV2 $T=837000 588120 0 0 $X=837000 $Y=587740
X3261 4590 873 1 2 INV2 $T=840100 578040 1 0 $X=840100 $Y=572620
X3262 4523 4594 1 2 INV2 $T=843820 699000 1 0 $X=843820 $Y=693580
X3263 916 4840 1 2 INV2 $T=879780 628440 0 0 $X=879780 $Y=628060
X3264 4875 4949 1 2 INV2 $T=897760 618360 0 0 $X=897760 $Y=617980
X3265 650 4875 1 2 INV2 $T=898380 719160 0 0 $X=898380 $Y=718780
X3266 5144 5159 1 2 INV2 $T=931860 638520 0 0 $X=931860 $Y=638140
X3267 5021 5171 1 2 INV2 $T=936820 608280 0 180 $X=934960 $Y=602860
X3268 5171 991 1 2 INV2 $T=939300 598200 1 0 $X=939300 $Y=592780
X3269 5240 1000 1 2 INV2 $T=947360 628440 1 180 $X=945500 $Y=628060
X3270 5159 5240 1 2 INV2 $T=947360 638520 1 180 $X=945500 $Y=638140
X3271 5266 5214 1 2 INV2 $T=951700 608280 1 0 $X=951700 $Y=602860
X3272 4650 5446 1 2 INV2 $T=987660 638520 1 0 $X=987660 $Y=633100
X3273 4650 1051 1 2 INV2 $T=989520 638520 1 0 $X=989520 $Y=633100
X3274 5422 5566 1 2 INV2 $T=1009360 588120 0 0 $X=1009360 $Y=587740
X3275 1841 1945 1 2 BUF2 $T=353400 668760 1 180 $X=350300 $Y=668380
X3276 462 3024 1 2 BUF2 $T=571640 578040 0 180 $X=568540 $Y=572620
X3277 3220 2920 1 2 BUF2 $T=584660 578040 1 180 $X=581560 $Y=577660
X3278 3192 3330 1 2 BUF2 $T=598920 578040 0 0 $X=598920 $Y=577660
X3279 620 650 1 2 BUF2 $T=654100 719160 0 0 $X=654100 $Y=718780
X3280 4148 3873 1 2 BUF2 $T=755780 638520 1 180 $X=752680 $Y=638140
X3281 4168 3859 1 2 BUF2 $T=758260 638520 0 0 $X=758260 $Y=638140
X3282 791 4164 1 2 BUF2 $T=767560 709080 0 0 $X=767560 $Y=708700
X3283 4253 4111 1 2 BUF2 $T=776860 648600 0 0 $X=776860 $Y=648220
X3284 4764 4910 1 2 BUF2 $T=889080 618360 0 0 $X=889080 $Y=617980
X3285 5034 5055 1 2 BUF2 $T=918220 658680 0 0 $X=918220 $Y=658300
X3286 5202 5219 1 2 BUF2 $T=941160 709080 0 0 $X=941160 $Y=708700
X3287 5894 5951 1 2 BUF2 $T=1075080 709080 0 0 $X=1075080 $Y=708700
X3288 16 1 18 19 2 17 ND3 $T=225680 719160 0 0 $X=225680 $Y=718780
X3289 1331 1 1284 1261 2 1296 ND3 $T=232500 699000 1 180 $X=230020 $Y=698620
X3290 31 1 1284 1340 2 1345 ND3 $T=240560 719160 1 180 $X=238080 $Y=718780
X3291 44 1 1387 1490 2 1404 ND3 $T=264120 557880 1 0 $X=264120 $Y=552460
X3292 1587 1 1469 1535 2 1579 ND3 $T=283340 557880 1 180 $X=280860 $Y=557500
X3293 211 1 210 166 2 2090 ND3 $T=396180 578040 0 180 $X=393700 $Y=572620
X3294 3369 1 3390 3450 2 2798 ND3 $T=623720 598200 0 0 $X=623720 $Y=597820
X3295 3457 1 2912 3429 2 2947 ND3 $T=628060 668760 0 180 $X=625580 $Y=663340
X3296 3494 1 3436 3514 2 613 ND3 $T=632400 688920 0 0 $X=632400 $Y=688540
X3297 593 1 3578 3597 2 3467 ND3 $T=649760 688920 1 180 $X=647280 $Y=688540
X3298 780 1 4223 792 2 783 ND3 $T=767560 719160 0 0 $X=767560 $Y=718780
X3299 4332 1 4449 4402 2 4454 ND3 $T=812820 678840 0 0 $X=812820 $Y=678460
X3300 4474 1 4472 841 2 3833 ND3 $T=819020 668760 0 180 $X=816540 $Y=663340
X3301 4480 1 4475 842 2 3874 ND3 $T=819640 668760 1 180 $X=817160 $Y=668380
X3302 4497 1 4489 846 2 3828 ND3 $T=821500 658680 1 180 $X=819020 $Y=658300
X3303 4699 1 4695 893 2 3939 ND3 $T=855600 668760 0 180 $X=853120 $Y=663340
X3304 4758 1 4748 906 2 3764 ND3 $T=864280 668760 1 180 $X=861800 $Y=668380
X3305 5030 1 5023 963 2 3865 ND3 $T=910780 567960 0 180 $X=908300 $Y=562540
X3306 5105 1 5097 976 2 3909 ND3 $T=925040 557880 0 180 $X=922560 $Y=552460
X3307 5108 1 978 977 2 3848 ND3 $T=925660 547800 0 180 $X=923180 $Y=542380
X3308 5112 1 5117 980 2 3825 ND3 $T=928140 588120 1 180 $X=925660 $Y=587740
X3309 5124 1 5118 981 2 3931 ND3 $T=928140 608280 1 180 $X=925660 $Y=607900
X3310 1284 1243 1291 2 1 ND2S $T=228160 699000 0 0 $X=228160 $Y=698620
X3311 1272 1331 1324 2 1 ND2S $T=233120 699000 0 0 $X=233120 $Y=698620
X3312 29 1343 10 2 1 ND2S $T=236220 537720 1 180 $X=234360 $Y=537340
X3313 28 1333 34 2 1 ND2S $T=240560 719160 0 0 $X=240560 $Y=718780
X3314 1404 1375 1413 2 1 ND2S $T=249860 557880 1 0 $X=249860 $Y=552460
X3315 1415 24 43 2 1 ND2S $T=251100 719160 0 0 $X=251100 $Y=718780
X3316 1462 1422 1469 2 1 ND2S $T=257920 537720 0 0 $X=257920 $Y=537340
X3317 1404 1467 1444 2 1 ND2S $T=259780 557880 1 0 $X=259780 $Y=552460
X3318 76 1550 1540 2 1 ND2S $T=275900 557880 1 0 $X=275900 $Y=552460
X3319 1497 1600 1562 2 1 ND2S $T=285200 588120 1 180 $X=283340 $Y=587740
X3320 1804 1741 1796 2 1 ND2S $T=319920 598200 0 0 $X=319920 $Y=597820
X3321 1930 1899 1935 2 1 ND2S $T=352160 678840 0 0 $X=352160 $Y=678460
X3322 1999 1936 2009 2 1 ND2S $T=363320 688920 1 0 $X=363320 $Y=683500
X3323 1974 1978 1973 2 1 ND2S $T=372000 547800 0 0 $X=372000 $Y=547420
X3324 1987 2230 2240 2 1 ND2S $T=404860 588120 1 0 $X=404860 $Y=582700
X3325 2070 2237 2232 2 1 ND2S $T=407340 578040 0 180 $X=405480 $Y=572620
X3326 2256 2300 1925 2 1 ND2S $T=419740 557880 1 180 $X=417880 $Y=557500
X3327 221 2303 2359 2 1 ND2S $T=423460 567960 1 0 $X=423460 $Y=562540
X3328 2331 2362 2287 2 1 ND2S $T=425320 567960 1 180 $X=423460 $Y=567580
X3329 2352 2365 2372 2 1 ND2S $T=426560 557880 0 0 $X=426560 $Y=557500
X3330 2355 2375 2362 2 1 ND2S $T=428420 578040 0 180 $X=426560 $Y=572620
X3331 2405 2412 2365 2 1 ND2S $T=434000 567960 1 0 $X=434000 $Y=562540
X3332 2411 2453 2286 2 1 ND2S $T=437720 547800 1 180 $X=435860 $Y=547420
X3333 247 2438 2439 2 1 ND2S $T=437720 537720 0 0 $X=437720 $Y=537340
X3334 2433 2439 2368 2 1 ND2S $T=439580 547800 1 180 $X=437720 $Y=547420
X3335 2427 2482 2453 2 1 ND2S $T=446400 547800 1 180 $X=444540 $Y=547420
X3336 369 366 368 2 1 ND2S $T=519560 537720 0 0 $X=519560 $Y=537340
X3337 2805 2932 2967 2 1 ND2S $T=530720 618360 1 0 $X=530720 $Y=612940
X3338 3069 3033 3073 2 1 ND2S $T=553040 628440 1 180 $X=551180 $Y=628060
X3339 3077 3061 3103 2 1 ND2S $T=560480 567960 1 180 $X=558620 $Y=567580
X3340 3106 3113 3122 2 1 ND2S $T=564200 557880 0 180 $X=562340 $Y=552460
X3341 3107 3234 3217 2 1 ND2S $T=585280 618360 1 180 $X=583420 $Y=617980
X3342 3172 3184 3262 2 1 ND2S $T=586520 598200 1 0 $X=586520 $Y=592780
X3343 3422 3397 587 2 1 ND2S $T=618760 688920 0 0 $X=618760 $Y=688540
X3344 3452 3426 2947 2 1 ND2S $T=625580 678840 1 0 $X=625580 $Y=673420
X3345 2798 3459 3303 2 1 ND2S $T=628060 608280 1 180 $X=626200 $Y=607900
X3346 2798 3485 3406 2 1 ND2S $T=629300 598200 1 180 $X=627440 $Y=597820
X3347 3434 3432 3510 2 1 ND2S $T=633020 699000 1 0 $X=633020 $Y=693580
X3348 3479 3489 2821 2 1 ND2S $T=633640 678840 0 0 $X=633640 $Y=678460
X3349 3543 3479 3494 2 1 ND2S $T=641700 688920 0 0 $X=641700 $Y=688540
X3350 3527 3480 3533 2 1 ND2S $T=647280 699000 0 0 $X=647280 $Y=698620
X3351 643 651 3528 2 1 ND2S $T=655960 557880 1 180 $X=654100 $Y=557500
X3352 3481 3706 3479 2 1 ND2S $T=668980 699000 1 180 $X=667120 $Y=698620
X3353 3726 3481 3610 2 1 ND2S $T=668980 699000 0 0 $X=668980 $Y=698620
X3354 3974 3590 3984 2 1 ND2S $T=721680 719160 1 0 $X=721680 $Y=713740
X3355 3706 3998 722 2 1 ND2S $T=722300 719160 0 0 $X=722300 $Y=718780
X3356 4005 728 3005 2 1 ND2S $T=732220 719160 1 0 $X=732220 $Y=713740
X3357 5516 5556 5542 2 1 ND2S $T=1006260 648600 1 180 $X=1004400 $Y=648220
X3358 1236 1235 1 1249 1260 1258 2 MOAI1S $T=220100 648600 1 0 $X=220100 $Y=643180
X3359 1244 1261 1 1244 1243 1238 2 MOAI1S $T=223820 699000 1 180 $X=220100 $Y=698620
X3360 1267 13 1 10 1245 1239 2 MOAI1S $T=224440 557880 0 180 $X=220720 $Y=552460
X3361 1242 1235 1 1249 1271 1250 2 MOAI1S $T=221960 658680 0 0 $X=221960 $Y=658300
X3362 1234 1272 1 1249 1281 1251 2 MOAI1S $T=223820 678840 0 0 $X=223820 $Y=678460
X3363 1241 1235 1 1282 1283 1301 2 MOAI1S $T=225060 628440 1 0 $X=225060 $Y=623020
X3364 1302 1259 1 1282 1286 1285 2 MOAI1S $T=231880 588120 1 180 $X=228160 $Y=587740
X3365 1237 1259 1 10 1279 1300 2 MOAI1S $T=229400 567960 0 0 $X=229400 $Y=567580
X3366 1319 1259 1 1282 1307 1303 2 MOAI1S $T=234980 598200 1 180 $X=231260 $Y=597820
X3367 1295 1259 1 1282 1298 1297 2 MOAI1S $T=231880 608280 1 0 $X=231880 $Y=602860
X3368 1314 1259 1 10 1328 1306 2 MOAI1S $T=233120 567960 1 0 $X=233120 $Y=562540
X3369 18 24 1 18 32 1384 2 MOAI1S $T=244280 719160 1 0 $X=244280 $Y=713740
X3370 1343 1380 1 1376 38 1262 2 MOAI1S $T=249240 537720 1 180 $X=245520 $Y=537340
X3371 1388 1387 1 1376 1375 1373 2 MOAI1S $T=249240 557880 0 180 $X=245520 $Y=552460
X3372 1343 41 1 1376 1422 1427 2 MOAI1S $T=249860 537720 0 0 $X=249860 $Y=537340
X3373 1388 44 1 1376 1445 1434 2 MOAI1S $T=252960 557880 0 0 $X=252960 $Y=557500
X3374 1460 47 1 1460 1456 1407 2 MOAI1S $T=259780 699000 1 180 $X=256060 $Y=698620
X3375 1460 51 1 1484 55 1487 2 MOAI1S $T=261020 699000 0 0 $X=261020 $Y=698620
X3376 1449 63 1 1449 1415 48 2 MOAI1S $T=269080 719160 1 180 $X=265360 $Y=718780
X3377 1502 1418 1 1483 1515 1486 2 MOAI1S $T=266600 638520 0 0 $X=266600 $Y=638140
X3378 70 66 1 70 67 1544 2 MOAI1S $T=271560 719160 1 0 $X=271560 $Y=713740
X3379 1525 1418 1 1483 1554 1546 2 MOAI1S $T=273420 638520 0 0 $X=273420 $Y=638140
X3380 70 75 1 70 1500 1569 2 MOAI1S $T=274040 709080 0 0 $X=274040 $Y=708700
X3381 1558 1565 1 1559 1529 1480 2 MOAI1S $T=279620 567960 1 180 $X=275900 $Y=567580
X3382 1558 1553 1 1560 1548 1503 2 MOAI1S $T=279620 578040 1 180 $X=275900 $Y=577660
X3383 1577 1566 1 1562 1561 1542 2 MOAI1S $T=279620 618360 1 180 $X=275900 $Y=617980
X3384 1484 80 1 1484 52 1563 2 MOAI1S $T=283340 699000 0 180 $X=279620 $Y=693580
X3385 1574 1566 1 1562 1596 1598 2 MOAI1S $T=280860 638520 1 0 $X=280860 $Y=633100
X3386 1568 1601 1 1560 1588 1505 2 MOAI1S $T=285820 578040 0 180 $X=282100 $Y=572620
X3387 1572 1558 1 1562 1602 1517 2 MOAI1S $T=282100 598200 1 0 $X=282100 $Y=592780
X3388 1558 1595 1 1559 1613 1476 2 MOAI1S $T=283960 567960 1 0 $X=283960 $Y=562540
X3389 1642 1566 1 1562 1627 1625 2 MOAI1S $T=293260 598200 0 180 $X=289540 $Y=592780
X3390 1652 1662 1 1652 90 1636 2 MOAI1S $T=296980 709080 1 180 $X=293260 $Y=708700
X3391 1652 1682 1 1652 106 1689 2 MOAI1S $T=299460 699000 1 0 $X=299460 $Y=693580
X3392 1695 1698 1 1695 91 1708 2 MOAI1S $T=303180 578040 0 0 $X=303180 $Y=577660
X3393 1484 103 1 1484 1723 1715 2 MOAI1S $T=310620 678840 1 180 $X=306900 $Y=678460
X3394 1652 1722 1 1652 116 1732 2 MOAI1S $T=306900 719160 1 0 $X=306900 $Y=713740
X3395 1734 1731 1 1649 1750 1753 2 MOAI1S $T=310620 588120 0 0 $X=310620 $Y=587740
X3396 1695 1751 1 1695 120 1710 2 MOAI1S $T=314340 678840 1 180 $X=310620 $Y=678460
X3397 1695 1764 1 1695 126 1717 2 MOAI1S $T=316820 578040 0 180 $X=313100 $Y=572620
X3398 1752 1756 1 1752 127 1779 2 MOAI1S $T=313100 709080 0 0 $X=313100 $Y=708700
X3399 1793 1418 1 1483 1767 1769 2 MOAI1S $T=321160 638520 1 180 $X=317440 $Y=638140
X3400 1752 1789 1 1752 68 1798 2 MOAI1S $T=318680 709080 1 0 $X=318680 $Y=703660
X3401 1783 1731 1 1649 1802 1792 2 MOAI1S $T=319920 588120 0 0 $X=319920 $Y=587740
X3402 1812 1817 1 1483 1827 1831 2 MOAI1S $T=324260 648600 0 0 $X=324260 $Y=648220
X3403 1794 1828 1 1794 118 1778 2 MOAI1S $T=327980 678840 1 180 $X=324260 $Y=678460
X3404 1810 1543 1 1849 1854 1760 2 MOAI1S $T=330460 678840 0 0 $X=330460 $Y=678460
X3405 1843 1418 1 1852 1837 1839 2 MOAI1S $T=331080 638520 1 0 $X=331080 $Y=633100
X3406 1860 1817 1 1852 1875 1872 2 MOAI1S $T=336040 648600 0 0 $X=336040 $Y=648220
X3407 1866 1731 1 1649 1879 1821 2 MOAI1S $T=337280 588120 0 0 $X=337280 $Y=587740
X3408 1885 153 1 1885 1883 1819 2 MOAI1S $T=343480 668760 1 180 $X=339760 $Y=668380
X3409 1895 1817 1 1852 1915 1921 2 MOAI1S $T=343480 628440 0 0 $X=343480 $Y=628060
X3410 1885 1922 1 1885 1835 1888 2 MOAI1S $T=347820 668760 1 180 $X=344100 $Y=668380
X3411 1903 1817 1 1852 1933 1909 2 MOAI1S $T=345960 648600 1 0 $X=345960 $Y=643180
X3412 1869 1835 1 1930 1935 1906 2 MOAI1S $T=345960 678840 0 0 $X=345960 $Y=678460
X3413 1942 1731 1 1649 1931 1924 2 MOAI1S $T=350920 588120 1 180 $X=347200 $Y=587740
X3414 1925 1593 1 88 1940 1927 2 MOAI1S $T=347200 608280 0 0 $X=347200 $Y=607900
X3415 1926 1817 1 1852 1918 1943 2 MOAI1S $T=347200 628440 0 0 $X=347200 $Y=628060
X3416 1914 1817 1 1852 1902 1944 2 MOAI1S $T=347200 638520 0 0 $X=347200 $Y=638140
X3417 1970 1731 1 1920 1959 1952 2 MOAI1S $T=356500 588120 1 180 $X=352780 $Y=587740
X3418 1794 1963 1 1794 174 1929 2 MOAI1S $T=354640 668760 0 0 $X=354640 $Y=668380
X3419 1841 1971 1 1841 1971 182 2 MOAI1S $T=358980 678840 0 0 $X=358980 $Y=678460
X3420 179 1998 1 179 177 2004 2 MOAI1S $T=362700 668760 1 0 $X=362700 $Y=663340
X3421 1987 2015 1 1920 2007 2002 2 MOAI1S $T=367660 588120 1 180 $X=363940 $Y=587740
X3422 1987 2035 1 1920 2042 2027 2 MOAI1S $T=368280 598200 1 0 $X=368280 $Y=592780
X3423 179 2037 1 179 187 2054 2 MOAI1S $T=369520 668760 1 0 $X=369520 $Y=663340
X3424 2014 1593 1 88 2028 2057 2 MOAI1S $T=370140 608280 0 0 $X=370140 $Y=607900
X3425 2128 1987 1 1920 2118 2114 2 MOAI1S $T=387500 588120 0 180 $X=383780 $Y=582700
X3426 2132 1987 1 1920 2147 2144 2 MOAI1S $T=387500 588120 1 0 $X=387500 $Y=582700
X3427 2130 2239 1 2207 2230 2223 2 MOAI1S $T=407340 588120 1 180 $X=403620 $Y=587740
X3428 2130 211 1 2248 2225 2267 2 MOAI1S $T=408580 578040 0 0 $X=408580 $Y=577660
X3429 3082 2708 1 3082 445 3140 2 MOAI1S $T=561720 709080 1 0 $X=561720 $Y=703660
X3430 3132 2971 1 3132 445 3134 2 MOAI1S $T=569780 709080 0 180 $X=566060 $Y=703660
X3431 3082 461 1 3082 3159 3128 2 MOAI1S $T=571640 719160 0 180 $X=567920 $Y=713740
X3432 3132 3183 1 3132 3159 3161 2 MOAI1S $T=574120 709080 0 180 $X=570400 $Y=703660
X3433 3132 477 1 3132 482 3210 2 MOAI1S $T=575980 719160 1 0 $X=575980 $Y=713740
X3434 3246 3255 1 3246 499 3257 2 MOAI1S $T=585900 709080 0 0 $X=585900 $Y=708700
X3435 432 495 1 432 499 3273 2 MOAI1S $T=585900 719160 1 0 $X=585900 $Y=713740
X3436 550 3358 1 550 544 540 2 MOAI1S $T=608840 719160 0 180 $X=605120 $Y=713740
X3437 3396 3395 1 3396 3395 2869 2 MOAI1S $T=617520 678840 0 180 $X=613800 $Y=673420
X3438 3368 2955 1 3368 3159 3340 2 MOAI1S $T=617520 709080 0 180 $X=613800 $Y=703660
X3439 3434 3421 1 3427 3421 3409 2 MOAI1S $T=621860 678840 1 180 $X=618140 $Y=678460
X3440 2912 3426 1 2912 3426 3357 2 MOAI1S $T=622480 668760 0 180 $X=618760 $Y=663340
X3441 3368 2914 1 3368 499 3387 2 MOAI1S $T=622480 709080 0 180 $X=618760 $Y=703660
X3442 3390 3428 1 3390 3428 3318 2 MOAI1S $T=623100 598200 1 180 $X=619380 $Y=597820
X3443 3430 3464 1 3430 3464 3175 2 MOAI1S $T=630540 598200 0 180 $X=626820 $Y=592780
X3444 3459 3450 1 3460 3430 3497 2 MOAI1S $T=627440 588120 0 0 $X=627440 $Y=587740
X3445 2947 593 1 2947 593 3487 2 MOAI1S $T=627440 678840 1 0 $X=627440 $Y=673420
X3446 3479 3342 1 3489 3498 3534 2 MOAI1S $T=629300 678840 0 0 $X=629300 $Y=678460
X3447 3450 3459 1 3450 3459 3511 2 MOAI1S $T=631160 598200 1 0 $X=631160 $Y=592780
X3448 3497 3485 1 3497 3485 3516 2 MOAI1S $T=631780 588120 0 0 $X=631780 $Y=587740
X3449 612 616 1 612 499 3473 2 MOAI1S $T=636740 719160 0 180 $X=633020 $Y=713740
X3450 3485 3497 1 3532 3557 632 2 MOAI1S $T=638600 578040 0 0 $X=638600 $Y=577660
X3451 3545 3546 1 3545 3546 3564 2 MOAI1S $T=640460 588120 1 0 $X=640460 $Y=582700
X3452 3590 3513 1 3573 3530 635 2 MOAI1S $T=648520 709080 0 180 $X=644800 $Y=703660
X3453 3553 3621 1 3553 3159 3596 2 MOAI1S $T=654720 678840 1 180 $X=651000 $Y=678460
X3454 3585 3652 1 3585 3613 3602 2 MOAI1S $T=660300 688920 1 180 $X=656580 $Y=688540
X3455 3630 3677 1 3630 3665 3648 2 MOAI1S $T=664020 638520 1 180 $X=660300 $Y=638140
X3456 3693 3635 1 3693 3665 3668 2 MOAI1S $T=668360 638520 1 180 $X=664640 $Y=638140
X3457 3694 3704 1 3694 3613 3664 2 MOAI1S $T=668360 668760 1 180 $X=664640 $Y=668380
X3458 3702 3683 1 3702 3613 3667 2 MOAI1S $T=669600 658680 1 180 $X=665880 $Y=658300
X3459 3595 3477 1 3595 3708 3634 2 MOAI1S $T=670840 578040 0 180 $X=667120 $Y=572620
X3460 3567 3715 1 3567 3665 3629 2 MOAI1S $T=670840 598200 0 180 $X=667120 $Y=592780
X3461 3713 3720 1 3713 3613 3684 2 MOAI1S $T=670840 688920 1 180 $X=667120 $Y=688540
X3462 3721 3418 1 3721 3708 3640 2 MOAI1S $T=672700 557880 0 180 $X=668980 $Y=552460
X3463 3702 3068 1 3702 3724 3669 2 MOAI1S $T=673940 658680 1 180 $X=670220 $Y=658300
X3464 3732 3739 1 3732 3613 3705 2 MOAI1S $T=675180 688920 1 180 $X=671460 $Y=688540
X3465 3721 3620 1 3721 667 3736 2 MOAI1S $T=677040 547800 0 180 $X=673320 $Y=542380
X3466 3741 3359 1 3741 3738 3637 2 MOAI1S $T=677040 567960 1 180 $X=673320 $Y=567580
X3467 3695 3756 1 3695 3665 3722 2 MOAI1S $T=677660 608280 0 180 $X=673940 $Y=602860
X3468 3694 3759 1 3694 3724 3744 2 MOAI1S $T=678280 658680 1 180 $X=674560 $Y=658300
X3469 3752 3763 1 3752 3665 3727 2 MOAI1S $T=678900 598200 0 180 $X=675180 $Y=592780
X3470 3630 3751 1 3630 3537 3767 2 MOAI1S $T=675180 638520 1 0 $X=675180 $Y=633100
X3471 3721 3772 1 3721 3738 3716 2 MOAI1S $T=680760 567960 0 180 $X=677040 $Y=562540
X3472 3693 3606 1 3693 3537 3765 2 MOAI1S $T=681380 638520 1 180 $X=677660 $Y=638140
X3473 3741 3775 1 3741 669 3731 2 MOAI1S $T=682000 557880 0 180 $X=678280 $Y=552460
X3474 3702 3778 1 3702 3768 3743 2 MOAI1S $T=682000 658680 1 180 $X=678280 $Y=658300
X3475 3694 3783 1 3694 3768 3746 2 MOAI1S $T=682620 668760 1 180 $X=678900 $Y=668380
X3476 3713 3135 1 3713 3768 3749 2 MOAI1S $T=683240 688920 1 180 $X=679520 $Y=688540
X3477 3695 3214 1 3695 3738 3712 2 MOAI1S $T=685100 618360 0 180 $X=681380 $Y=612940
X3478 3776 3521 1 3776 679 3717 2 MOAI1S $T=685720 578040 1 180 $X=682000 $Y=577660
X3479 3792 3623 1 3792 679 3718 2 MOAI1S $T=686340 588120 0 180 $X=682620 $Y=582700
X3480 3732 3807 1 3732 3768 3766 2 MOAI1S $T=687580 688920 1 180 $X=683860 $Y=688540
X3481 3752 3711 1 3752 3738 3785 2 MOAI1S $T=688820 618360 0 180 $X=685100 $Y=612940
X3482 3741 684 1 3741 667 3816 2 MOAI1S $T=686340 547800 0 0 $X=686340 $Y=547420
X3483 685 688 1 685 667 690 2 MOAI1S $T=688200 537720 0 0 $X=688200 $Y=537340
X3484 3847 3836 1 3847 3738 3840 2 MOAI1S $T=696880 578040 0 180 $X=693160 $Y=572620
X3485 3858 3867 1 3858 669 3829 2 MOAI1S $T=698740 557880 0 180 $X=695020 $Y=552460
X3486 3858 3697 1 3858 698 3839 2 MOAI1S $T=695640 557880 0 0 $X=695640 $Y=557500
X3487 3824 3901 1 3824 703 3884 2 MOAI1S $T=706180 668760 1 180 $X=702460 $Y=668380
X3488 3858 3470 1 3858 701 3882 2 MOAI1S $T=706800 547800 1 180 $X=703080 $Y=547420
X3489 3862 3302 1 3862 3658 3879 2 MOAI1S $T=707420 618360 0 180 $X=703700 $Y=612940
X3490 3811 3655 1 3811 3658 3896 2 MOAI1S $T=709280 638520 0 180 $X=705560 $Y=633100
X3491 3843 3222 1 3843 3658 3891 2 MOAI1S $T=709280 658680 1 180 $X=705560 $Y=658300
X3492 3897 3117 1 3897 703 3871 2 MOAI1S $T=709900 688920 0 180 $X=706180 $Y=683500
X3493 3890 3911 1 3890 3658 3934 2 MOAI1S $T=709280 638520 1 0 $X=709280 $Y=633100
X3494 3916 3685 1 3916 669 3940 2 MOAI1S $T=710520 557880 1 0 $X=710520 $Y=552460
X3495 3916 3920 1 3916 701 3932 2 MOAI1S $T=710520 567960 0 0 $X=710520 $Y=567580
X3496 3885 3570 1 3885 701 3937 2 MOAI1S $T=711140 618360 1 0 $X=711140 $Y=612940
X3497 3918 3035 1 3918 703 3922 2 MOAI1S $T=714860 709080 0 180 $X=711140 $Y=703660
X3498 3005 727 1 3005 3998 4035 2 MOAI1S $T=729120 719160 0 0 $X=729120 $Y=718780
X3499 4129 771 1 720 4122 4089 2 MOAI1S $T=752060 719160 1 180 $X=748340 $Y=718780
X3500 4479 4450 1 4479 4476 4469 2 MOAI1S $T=821500 709080 0 180 $X=817780 $Y=703660
X3501 4486 4495 1 4486 4476 4468 2 MOAI1S $T=822740 699000 0 180 $X=819020 $Y=693580
X3502 4494 3453 1 4494 4476 4465 2 MOAI1S $T=823980 688920 1 180 $X=820260 $Y=688540
X3503 4508 4519 1 4508 4476 4482 2 MOAI1S $T=827080 648600 0 180 $X=823360 $Y=643180
X3504 4528 3491 1 4528 4476 4453 2 MOAI1S $T=829560 678840 0 180 $X=825840 $Y=673420
X3505 4562 3548 1 4508 4521 4448 2 MOAI1S $T=830800 648600 1 180 $X=827080 $Y=648220
X3506 4556 4511 1 4556 4568 4563 2 MOAI1S $T=830180 699000 0 0 $X=830180 $Y=698620
X3507 4508 874 1 4508 4599 4551 2 MOAI1S $T=840720 628440 1 180 $X=837000 $Y=628060
X3508 4550 4607 1 4610 4521 4620 2 MOAI1S $T=838240 648600 0 0 $X=838240 $Y=648220
X3509 4486 4626 1 4486 4521 4605 2 MOAI1S $T=843820 699000 0 180 $X=840100 $Y=693580
X3510 4550 3566 1 4550 4599 4653 2 MOAI1S $T=840720 628440 0 0 $X=840720 $Y=628060
X3511 4528 4623 1 4528 4521 4635 2 MOAI1S $T=841340 668760 0 0 $X=841340 $Y=668380
X3512 4544 4661 1 4544 4521 4638 2 MOAI1S $T=849400 709080 0 180 $X=845680 $Y=703660
X3513 4494 4543 1 4494 4521 4631 2 MOAI1S $T=850020 688920 0 180 $X=846300 $Y=683500
X3514 4610 4665 1 4610 4654 4634 2 MOAI1S $T=850640 648600 1 180 $X=846920 $Y=648220
X3515 4660 4715 1 4660 4719 4732 2 MOAI1S $T=856220 658680 0 0 $X=856220 $Y=658300
X3516 4486 4717 1 4725 4719 4740 2 MOAI1S $T=856220 699000 1 0 $X=856220 $Y=693580
X3517 4727 4737 1 4727 4654 4643 2 MOAI1S $T=861180 638520 1 180 $X=857460 $Y=638140
X3518 4544 4722 1 4733 4719 4662 2 MOAI1S $T=862420 709080 1 180 $X=858700 $Y=708700
X3519 4731 4639 1 4731 4745 4746 2 MOAI1S $T=859320 628440 0 0 $X=859320 $Y=628060
X3520 4673 4749 1 4744 4719 4741 2 MOAI1S $T=864280 678840 0 180 $X=860560 $Y=673420
X3521 4727 4747 1 4727 910 4770 2 MOAI1S $T=862420 638520 0 0 $X=862420 $Y=638140
X3522 4701 4768 1 4701 4719 4753 2 MOAI1S $T=867380 688920 0 180 $X=863660 $Y=683500
X3523 4725 4788 1 4725 916 4769 2 MOAI1S $T=871720 688920 1 180 $X=868000 $Y=688540
X3524 4701 4804 1 4701 916 4792 2 MOAI1S $T=874820 688920 0 180 $X=871100 $Y=683500
X3525 4799 4671 1 4799 4714 4789 2 MOAI1S $T=875440 628440 0 180 $X=871720 $Y=623020
X3526 4744 4812 1 4744 916 4830 2 MOAI1S $T=874200 678840 1 0 $X=874200 $Y=673420
X3527 4578 4836 1 4578 924 4765 2 MOAI1S $T=880400 608280 1 180 $X=876680 $Y=607900
X3528 4822 4825 1 4822 916 4835 2 MOAI1S $T=876680 648600 1 0 $X=876680 $Y=643180
X3529 4733 4837 1 4733 916 4816 2 MOAI1S $T=880400 709080 1 180 $X=876680 $Y=708700
X3530 4831 4849 1 4831 925 4814 2 MOAI1S $T=882260 598200 0 180 $X=878540 $Y=592780
X3531 4856 4865 1 4856 924 4839 2 MOAI1S $T=884740 608280 1 180 $X=881020 $Y=607900
X3532 4733 4881 1 4733 930 4826 2 MOAI1S $T=886600 709080 1 180 $X=882880 $Y=708700
X3533 4725 4890 1 4725 4900 4907 2 MOAI1S $T=886600 699000 1 0 $X=886600 $Y=693580
X3534 4888 4904 1 4888 925 4860 2 MOAI1S $T=890940 608280 0 180 $X=887220 $Y=602860
X3535 4660 4906 1 4660 4903 4921 2 MOAI1S $T=889080 658680 0 0 $X=889080 $Y=658300
X3536 4744 4895 1 4744 4900 4874 2 MOAI1S $T=892800 668760 1 180 $X=889080 $Y=668380
X3537 4672 4926 1 4672 4903 4939 2 MOAI1S $T=892800 658680 0 0 $X=892800 $Y=658300
X3538 4888 4936 1 4888 4944 4945 2 MOAI1S $T=894660 578040 0 0 $X=894660 $Y=577660
X3539 4917 945 1 4917 4714 4924 2 MOAI1S $T=899620 557880 0 180 $X=895900 $Y=552460
X3540 4959 949 1 4959 947 4891 2 MOAI1S $T=902720 537720 1 180 $X=899000 $Y=537340
X3541 4959 950 1 4959 4944 4901 2 MOAI1S $T=902720 578040 1 180 $X=899000 $Y=577660
X3542 4917 4933 1 4917 4967 4892 2 MOAI1S $T=900240 557880 0 0 $X=900240 $Y=557500
X3543 4831 957 1 4831 4967 4918 2 MOAI1S $T=905200 578040 0 180 $X=901480 $Y=572620
X3544 4959 5022 1 4959 4599 966 2 MOAI1S $T=910160 537720 0 0 $X=910160 $Y=537340
X3545 4925 4983 1 4925 4944 4986 2 MOAI1S $T=913880 578040 0 180 $X=910160 $Y=572620
X3546 5037 5044 1 5037 4599 5032 2 MOAI1S $T=915120 547800 1 180 $X=911400 $Y=547420
X3547 5037 5047 1 5037 4967 5026 2 MOAI1S $T=915120 567960 0 180 $X=911400 $Y=562540
X3548 5037 5057 1 5037 4714 5066 2 MOAI1S $T=915120 567960 1 0 $X=915120 $Y=562540
X3549 4943 5075 1 4943 4944 5045 2 MOAI1S $T=921320 578040 1 180 $X=917600 $Y=577660
X3550 5073 972 1 5073 4599 5099 2 MOAI1S $T=919460 547800 1 0 $X=919460 $Y=542380
X3551 5073 5062 1 5073 4967 5094 2 MOAI1S $T=927520 567960 0 180 $X=923800 $Y=562540
X3552 4658 5130 1 4658 5100 5109 2 MOAI1S $T=933720 578040 0 180 $X=930000 $Y=572620
X3553 5151 5154 1 879 985 5120 2 MOAI1S $T=934960 598200 0 180 $X=931240 $Y=592780
X3554 5149 5162 1 5149 987 5114 2 MOAI1S $T=935580 547800 0 180 $X=931860 $Y=542380
X3555 5073 988 1 5073 5167 5169 2 MOAI1S $T=932480 547800 0 0 $X=932480 $Y=547420
X3556 5149 5195 1 5149 4967 5208 2 MOAI1S $T=938680 567960 1 0 $X=938680 $Y=562540
X3557 5194 995 1 5194 987 5213 2 MOAI1S $T=939300 547800 1 0 $X=939300 $Y=542380
X3558 5149 5200 1 5149 5167 5215 2 MOAI1S $T=940540 557880 1 0 $X=940540 $Y=552460
X3559 5151 5209 1 5151 5100 5248 2 MOAI1S $T=942400 588120 1 0 $X=942400 $Y=582700
X3560 5194 5234 1 5194 5167 5268 2 MOAI1S $T=945500 557880 1 0 $X=945500 $Y=552460
X3561 5207 5235 1 5207 985 5252 2 MOAI1S $T=945500 598200 1 0 $X=945500 $Y=592780
X3562 5194 5246 1 5194 4967 5259 2 MOAI1S $T=947360 567960 0 0 $X=947360 $Y=567580
X3563 5278 1006 1 5278 1011 5267 2 MOAI1S $T=952940 547800 1 0 $X=952940 $Y=542380
X3564 5278 1013 1 5278 5303 5307 2 MOAI1S $T=956660 547800 1 0 $X=956660 $Y=542380
X3565 5278 5297 1 5278 5167 5314 2 MOAI1S $T=959760 557880 0 0 $X=959760 $Y=557500
X3566 5308 1018 1 5308 1011 5318 2 MOAI1S $T=960380 547800 1 0 $X=960380 $Y=542380
X3567 5308 5319 1 5308 5167 5330 2 MOAI1S $T=962240 567960 1 0 $X=962240 $Y=562540
X3568 5308 1019 1 5308 5303 5334 2 MOAI1S $T=964100 547800 1 0 $X=964100 $Y=542380
X3569 5374 5389 1 5374 5375 5373 2 MOAI1S $T=981460 658680 0 180 $X=977740 $Y=653260
X3570 5374 5390 1 5374 4900 5344 2 MOAI1S $T=981460 668760 1 180 $X=977740 $Y=668380
X3571 5379 5356 1 5379 4900 5352 2 MOAI1S $T=981460 678840 1 180 $X=977740 $Y=678460
X3572 5379 5376 1 5379 5375 5329 2 MOAI1S $T=982700 658680 1 180 $X=978980 $Y=658300
X3573 5407 1040 1 5407 1033 5343 2 MOAI1S $T=985800 547800 1 180 $X=982080 $Y=547420
X3574 5408 5415 1 5408 5100 5366 2 MOAI1S $T=985800 588120 0 180 $X=982080 $Y=582700
X3575 5414 5357 1 5414 4903 5353 2 MOAI1S $T=987040 709080 0 180 $X=983320 $Y=703660
X3576 5443 5437 1 5407 5358 5339 2 MOAI1S $T=988900 567960 1 180 $X=985180 $Y=567580
X3577 1028 5392 1 1028 974 5378 2 MOAI1S $T=990140 557880 0 180 $X=986420 $Y=552460
X3578 5368 5461 1 5368 1055 5434 2 MOAI1S $T=992620 688920 1 180 $X=988900 $Y=688540
X3579 5408 1067 1 5408 974 5395 2 MOAI1S $T=993860 557880 0 180 $X=990140 $Y=552460
X3580 5407 1064 1 5407 1069 1071 2 MOAI1S $T=991380 537720 0 0 $X=991380 $Y=537340
X3581 5448 1070 1 5448 1033 1062 2 MOAI1S $T=995100 547800 0 180 $X=991380 $Y=542380
X3582 5414 5479 1 5414 1055 5463 2 MOAI1S $T=995100 709080 0 180 $X=991380 $Y=703660
X3583 5494 5505 1 5494 5358 5480 2 MOAI1S $T=999440 608280 1 180 $X=995720 $Y=607900
X3584 5469 5513 1 5469 1055 5528 2 MOAI1S $T=998820 678840 0 0 $X=998820 $Y=678460
X3585 5522 5529 1 5522 5358 5495 2 MOAI1S $T=1003780 608280 1 180 $X=1000060 $Y=607900
X3586 5350 5531 1 5350 5519 5510 2 MOAI1S $T=1003780 638520 0 180 $X=1000060 $Y=633100
X3587 5368 5532 1 5368 1081 5507 2 MOAI1S $T=1004400 699000 0 180 $X=1000680 $Y=693580
X3588 5443 5436 1 5443 974 5493 2 MOAI1S $T=1005640 557880 1 180 $X=1001920 $Y=557500
X3589 5469 5459 1 5469 5519 5501 2 MOAI1S $T=1006880 678840 1 180 $X=1003160 $Y=678460
X3590 5442 5557 1 5442 1081 5508 2 MOAI1S $T=1007500 709080 1 180 $X=1003780 $Y=708700
X3591 5547 5559 1 5547 5100 5536 2 MOAI1S $T=1008120 578040 0 180 $X=1004400 $Y=572620
X3592 1072 5549 1 1072 974 5564 2 MOAI1S $T=1005020 547800 0 0 $X=1005020 $Y=547420
X3593 5539 5567 1 5539 985 5551 2 MOAI1S $T=1009360 588120 1 180 $X=1005640 $Y=587740
X3594 5385 5571 1 5385 5519 5553 2 MOAI1S $T=1009980 668760 1 180 $X=1006260 $Y=668380
X3595 5581 5466 1 5466 5519 5552 2 MOAI1S $T=1010600 648600 1 180 $X=1006880 $Y=648220
X3596 5412 5576 1 5412 5519 5596 2 MOAI1S $T=1008740 638520 1 0 $X=1008740 $Y=633100
X3597 1075 5586 1 1075 1086 1085 2 MOAI1S $T=1012460 719160 1 180 $X=1008740 $Y=718780
X3598 5448 5580 1 5448 1069 1092 2 MOAI1S $T=1009980 537720 0 0 $X=1009980 $Y=537340
X3599 5582 5591 1 5582 5519 5563 2 MOAI1S $T=1013700 688920 0 180 $X=1009980 $Y=683500
X3600 1091 5604 1 1091 1090 5587 2 MOAI1S $T=1015560 557880 0 180 $X=1011840 $Y=552460
X3601 5597 5603 1 5597 5574 5618 2 MOAI1S $T=1013700 547800 0 0 $X=1013700 $Y=547420
X3602 5597 1094 1 5597 1069 1095 2 MOAI1S $T=1014320 537720 0 0 $X=1014320 $Y=537340
X3603 5619 5629 1 5619 5100 5607 2 MOAI1S $T=1018660 578040 0 180 $X=1014940 $Y=572620
X3604 5625 5630 1 5625 5623 5593 2 MOAI1S $T=1019280 638520 0 180 $X=1015560 $Y=633100
X3605 5578 5631 1 5578 5623 5613 2 MOAI1S $T=1019280 678840 1 180 $X=1015560 $Y=678460
X3606 1091 1096 1 1091 5574 5621 2 MOAI1S $T=1019900 557880 0 180 $X=1016180 $Y=552460
X3607 5612 5626 1 5612 5623 5639 2 MOAI1S $T=1016180 648600 0 0 $X=1016180 $Y=648220
X3608 5610 5635 1 5610 1086 5617 2 MOAI1S $T=1019900 709080 1 180 $X=1016180 $Y=708700
X3609 5638 5643 1 5638 1090 5653 2 MOAI1S $T=1019280 557880 0 0 $X=1019280 $Y=557500
X3610 5590 5645 1 5590 5623 5656 2 MOAI1S $T=1019280 678840 0 0 $X=1019280 $Y=678460
X3611 5608 5620 1 5608 5623 5595 2 MOAI1S $T=1024240 628440 1 180 $X=1020520 $Y=628060
X3612 5605 5647 1 5605 1086 5662 2 MOAI1S $T=1020520 699000 1 0 $X=1020520 $Y=693580
X3613 5579 5660 1 5579 5623 5676 2 MOAI1S $T=1022380 658680 0 0 $X=1022380 $Y=658300
X3614 5625 5664 1 5625 5674 5668 2 MOAI1S $T=1028580 628440 1 180 $X=1024860 $Y=628060
X3615 5578 5677 1 5578 5674 5696 2 MOAI1S $T=1025480 678840 0 0 $X=1025480 $Y=678460
X3616 1109 5697 1 1109 5637 5729 2 MOAI1S $T=1029200 537720 0 0 $X=1029200 $Y=537340
X3617 1110 1112 1 1110 5637 5707 2 MOAI1S $T=1029200 547800 0 0 $X=1029200 $Y=547420
X3618 1110 1113 1 1110 5705 5709 2 MOAI1S $T=1029200 557880 0 0 $X=1029200 $Y=557500
X3619 5605 5699 1 5605 1111 5712 2 MOAI1S $T=1029200 699000 1 0 $X=1029200 $Y=693580
X3620 5612 5706 1 5612 5674 5734 2 MOAI1S $T=1031060 648600 0 0 $X=1031060 $Y=648220
X3621 5579 5710 1 5579 5674 5722 2 MOAI1S $T=1032300 658680 0 0 $X=1032300 $Y=658300
X3622 5714 5608 1 5608 5674 5718 2 MOAI1S $T=1032920 628440 0 0 $X=1032920 $Y=628060
X3623 5590 5723 1 5590 5674 5711 2 MOAI1S $T=1036640 678840 0 180 $X=1032920 $Y=673420
X3624 1109 5728 1 1109 5705 5740 2 MOAI1S $T=1035400 557880 0 0 $X=1035400 $Y=557500
X3625 5610 5733 1 5610 1111 5713 2 MOAI1S $T=1040980 709080 0 180 $X=1037260 $Y=703660
X3626 24 2 1272 1321 1 NR2 $T=233120 709080 1 0 $X=233120 $Y=703660
X3627 23 2 25 19 1 NR2 $T=233120 719160 0 0 $X=233120 $Y=718780
X3628 30 2 1345 1350 1 NR2 $T=238700 719160 1 0 $X=238700 $Y=713740
X3629 31 2 34 33 1 NR2 $T=244280 719160 1 180 $X=242420 $Y=718780
X3630 1414 2 1377 1397 1 NR2 $T=251100 588120 1 180 $X=249240 $Y=587740
X3631 1398 2 1389 1408 1 NR2 $T=249240 598200 1 0 $X=249240 $Y=592780
X3632 1399 2 1385 1410 1 NR2 $T=249240 628440 0 0 $X=249240 $Y=628060
X3633 1399 2 1391 1397 1 NR2 $T=249240 648600 1 0 $X=249240 $Y=643180
X3634 1399 2 1365 1398 1 NR2 $T=249240 658680 1 0 $X=249240 $Y=653260
X3635 42 2 1400 1393 1 NR2 $T=251100 699000 0 180 $X=249240 $Y=693580
X3636 1409 2 1249 1396 1 NR2 $T=251100 719160 0 180 $X=249240 $Y=713740
X3637 1424 2 1431 1414 1 NR2 $T=252960 598200 1 180 $X=251100 $Y=597820
X3638 1424 2 1416 1397 1 NR2 $T=252960 638520 0 180 $X=251100 $Y=633100
X3639 1414 2 1439 1410 1 NR2 $T=252960 588120 1 0 $X=252960 $Y=582700
X3640 1421 2 1432 1437 1 NR2 $T=252960 658680 1 0 $X=252960 $Y=653260
X3641 1425 2 1446 1441 1 NR2 $T=254200 648600 1 0 $X=254200 $Y=643180
X3642 1410 2 1471 1397 1 NR2 $T=256680 598200 1 180 $X=254820 $Y=597820
X3643 1437 2 1433 1455 1 NR2 $T=254820 678840 1 0 $X=254820 $Y=673420
X3644 1410 2 1450 1408 1 NR2 $T=255440 588120 1 0 $X=255440 $Y=582700
X3645 1410 2 1436 1398 1 NR2 $T=256680 608280 0 0 $X=256680 $Y=607900
X3646 1397 2 1458 1398 1 NR2 $T=256680 628440 0 0 $X=256680 $Y=628060
X3647 1425 2 1440 1437 1 NR2 $T=256680 638520 1 0 $X=256680 $Y=633100
X3648 1424 2 1470 1398 1 NR2 $T=256680 648600 1 0 $X=256680 $Y=643180
X3649 1421 2 1447 1441 1 NR2 $T=258540 658680 0 180 $X=256680 $Y=653260
X3650 1464 2 1472 1437 1 NR2 $T=258540 668760 0 180 $X=256680 $Y=663340
X3651 1425 2 1448 1454 1 NR2 $T=258540 668760 1 180 $X=256680 $Y=668380
X3652 1441 2 1426 1464 1 NR2 $T=256680 678840 0 0 $X=256680 $Y=678460
X3653 1428 2 1459 1464 1 NR2 $T=256680 699000 1 0 $X=256680 $Y=693580
X3654 1425 2 1475 52 1 NR2 $T=257920 678840 1 0 $X=257920 $Y=673420
X3655 1399 2 1466 1437 1 NR2 $T=260400 608280 1 180 $X=258540 $Y=607900
X3656 1421 2 1474 1454 1 NR2 $T=258540 668760 0 0 $X=258540 $Y=668380
X3657 1456 2 1457 1399 1 NR2 $T=260400 688920 0 180 $X=258540 $Y=683500
X3658 1399 2 1473 1443 1 NR2 $T=259780 628440 0 0 $X=259780 $Y=628060
X3659 1441 2 1477 1455 1 NR2 $T=259780 699000 1 0 $X=259780 $Y=693580
X3660 1456 2 1481 1425 1 NR2 $T=263500 688920 1 180 $X=261640 $Y=688540
X3661 1424 2 1493 1408 1 NR2 $T=265980 608280 0 180 $X=264120 $Y=602860
X3662 1424 2 1468 1410 1 NR2 $T=265980 618360 1 180 $X=264120 $Y=617980
X3663 1500 2 1495 1464 1 NR2 $T=266600 699000 0 180 $X=264740 $Y=693580
X3664 1443 2 1498 1398 1 NR2 $T=265360 608280 0 0 $X=265360 $Y=607900
X3665 1441 2 1516 1393 1 NR2 $T=269080 688920 0 0 $X=269080 $Y=688540
X3666 1528 2 1537 1535 1 NR2 $T=272180 567960 1 0 $X=272180 $Y=562540
X3667 1428 2 1538 1455 1 NR2 $T=272180 688920 0 0 $X=272180 $Y=688540
X3668 1550 2 1404 1535 1 NR2 $T=275900 557880 0 180 $X=274040 $Y=552460
X3669 73 2 1553 1490 1 NR2 $T=274040 578040 1 0 $X=274040 $Y=572620
X3670 1556 2 1573 79 1 NR2 $T=277760 688920 0 0 $X=277760 $Y=688540
X3671 1421 2 1555 52 1 NR2 $T=280860 658680 1 180 $X=279000 $Y=658300
X3672 1540 2 1595 1535 1 NR2 $T=281480 567960 1 0 $X=281480 $Y=562540
X3673 1428 2 1594 1393 1 NR2 $T=283960 699000 1 0 $X=283960 $Y=693580
X3674 1454 2 1615 1455 1 NR2 $T=290160 668760 1 180 $X=288300 $Y=668380
X3675 1454 2 1639 1629 1 NR2 $T=290160 668760 1 0 $X=290160 $Y=663340
X3676 1501 2 1630 1543 1 NR2 $T=293880 668760 1 180 $X=292020 $Y=668380
X3677 1651 2 1640 94 1 NR2 $T=293880 678840 1 180 $X=292020 $Y=678460
X3678 1501 2 1667 1656 1 NR2 $T=293880 668760 1 0 $X=293880 $Y=663340
X3679 1651 2 1647 1455 1 NR2 $T=297600 668760 1 180 $X=295740 $Y=668380
X3680 1501 2 1643 1629 1 NR2 $T=299460 668760 0 180 $X=297600 $Y=663340
X3681 1692 2 1686 1464 1 NR2 $T=300700 638520 1 180 $X=298840 $Y=638140
X3682 1501 2 1671 1464 1 NR2 $T=300700 658680 0 180 $X=298840 $Y=653260
X3683 1651 2 1678 1629 1 NR2 $T=301940 668760 0 180 $X=300080 $Y=663340
X3684 1692 2 1694 1712 1 NR2 $T=304420 618360 0 0 $X=304420 $Y=617980
X3685 1702 2 1696 1701 1 NR2 $T=306280 628440 1 180 $X=304420 $Y=628060
X3686 1702 2 1693 1721 1 NR2 $T=305660 638520 0 0 $X=305660 $Y=638140
X3687 1702 2 1724 1712 1 NR2 $T=306280 618360 1 0 $X=306280 $Y=612940
X3688 1692 2 1628 1721 1 NR2 $T=309380 638520 1 180 $X=307520 $Y=638140
X3689 1692 2 1746 1758 1 NR2 $T=311860 628440 1 0 $X=311860 $Y=623020
X3690 1721 2 1754 1701 1 NR2 $T=314960 618360 1 0 $X=314960 $Y=612940
X3691 1702 2 1773 1758 1 NR2 $T=314960 618360 0 0 $X=314960 $Y=617980
X3692 1701 2 1832 1712 1 NR2 $T=332940 608280 0 0 $X=332940 $Y=607900
X3693 1701 2 1913 1758 1 NR2 $T=343480 618360 1 0 $X=343480 $Y=612940
X3694 1758 2 1928 1712 1 NR2 $T=349060 618360 0 180 $X=347200 $Y=612940
X3695 162 2 1910 1936 1 NR2 $T=350300 719160 0 180 $X=348440 $Y=713740
X3696 167 2 1947 1936 1 NR2 $T=352780 719160 0 180 $X=350920 $Y=713740
X3697 162 2 168 1951 1 NR2 $T=350920 719160 0 0 $X=350920 $Y=718780
X3698 183 2 1938 1936 1 NR2 $T=364560 709080 1 180 $X=362700 $Y=708700
X3699 183 2 2011 1951 1 NR2 $T=364560 709080 0 0 $X=364560 $Y=708700
X3700 167 2 2024 1951 1 NR2 $T=368900 709080 1 180 $X=367040 $Y=708700
X3701 188 2 2021 1951 1 NR2 $T=370140 688920 1 180 $X=368280 $Y=688540
X3702 198 2 2080 192 1 NR2 $T=377580 699000 0 180 $X=375720 $Y=693580
X3703 188 2 2086 192 1 NR2 $T=380060 719160 0 180 $X=378200 $Y=713740
X3704 188 2 2069 191 1 NR2 $T=380680 719160 1 0 $X=380680 $Y=713740
X3705 198 2 2092 191 1 NR2 $T=382540 699000 1 0 $X=382540 $Y=693580
X3706 199 2 2105 197 1 NR2 $T=384400 709080 1 180 $X=382540 $Y=708700
X3707 199 2 2102 204 1 NR2 $T=384400 719160 1 0 $X=384400 $Y=713740
X3708 2143 2 2141 191 1 NR2 $T=390600 678840 1 180 $X=388740 $Y=678460
X3709 207 2 2125 2096 1 NR2 $T=389980 709080 0 0 $X=389980 $Y=708700
X3710 2169 2 2168 2096 1 NR2 $T=393080 699000 1 180 $X=391220 $Y=698620
X3711 2169 2 2160 203 1 NR2 $T=393700 709080 1 180 $X=391840 $Y=708700
X3712 2181 2 2175 203 1 NR2 $T=395560 699000 1 180 $X=393700 $Y=698620
X3713 2169 2 2166 208 1 NR2 $T=394940 709080 0 0 $X=394940 $Y=708700
X3714 2181 2 2187 212 1 NR2 $T=396180 699000 0 0 $X=396180 $Y=698620
X3715 207 2 2178 2121 1 NR2 $T=398660 688920 0 180 $X=396800 $Y=683500
X3716 2196 2 2180 212 1 NR2 $T=399280 678840 1 180 $X=397420 $Y=678460
X3717 2181 2 2235 213 1 NR2 $T=398660 699000 1 0 $X=398660 $Y=693580
X3718 2169 2 2200 212 1 NR2 $T=398660 709080 0 0 $X=398660 $Y=708700
X3719 207 2 2201 212 1 NR2 $T=398660 719160 1 0 $X=398660 $Y=713740
X3720 207 2 2184 213 1 NR2 $T=402380 719160 0 180 $X=400520 $Y=713740
X3721 214 2 215 216 1 NR2 $T=402380 537720 0 0 $X=402380 $Y=537340
X3722 2169 2 2241 213 1 NR2 $T=406100 719160 0 180 $X=404240 $Y=713740
X3723 2266 2 2246 2154 1 NR2 $T=409200 668760 0 180 $X=407340 $Y=663340
X3724 2181 2 2231 208 1 NR2 $T=409200 699000 1 180 $X=407340 $Y=698620
X3725 2259 2 2222 208 1 NR2 $T=410440 678840 1 180 $X=408580 $Y=678460
X3726 2259 2 2249 213 1 NR2 $T=412300 678840 1 180 $X=410440 $Y=678460
X3727 2265 2 2281 222 1 NR2 $T=412300 699000 1 180 $X=410440 $Y=698620
X3728 2265 2 2276 2277 1 NR2 $T=411060 699000 1 0 $X=411060 $Y=693580
X3729 2254 2 2293 2277 1 NR2 $T=414780 709080 0 180 $X=412920 $Y=703660
X3730 231 2 2289 2277 1 NR2 $T=414780 719160 1 180 $X=412920 $Y=718780
X3731 2294 2 2279 2277 1 NR2 $T=416020 688920 0 180 $X=414160 $Y=683500
X3732 214 2 2299 232 1 NR2 $T=415400 547800 1 0 $X=415400 $Y=542380
X3733 216 2 2307 232 1 NR2 $T=416020 557880 0 0 $X=416020 $Y=557500
X3734 2259 2 2295 229 1 NR2 $T=416640 678840 1 0 $X=416640 $Y=673420
X3735 2294 2 2296 229 1 NR2 $T=416640 688920 1 0 $X=416640 $Y=683500
X3736 2265 2 2337 236 1 NR2 $T=421600 709080 1 0 $X=421600 $Y=703660
X3737 2259 2 2320 2277 1 NR2 $T=422220 678840 1 0 $X=422220 $Y=673420
X3738 2294 2 2343 236 1 NR2 $T=422840 688920 1 0 $X=422840 $Y=683500
X3739 2294 2 2364 222 1 NR2 $T=423460 688920 0 0 $X=423460 $Y=688540
X3740 2254 2 2344 236 1 NR2 $T=425320 709080 0 180 $X=423460 $Y=703660
X3741 2266 2 2335 229 1 NR2 $T=425940 668760 0 180 $X=424080 $Y=663340
X3742 2181 2 2371 2342 1 NR2 $T=424700 699000 1 0 $X=424700 $Y=693580
X3743 231 2 2340 236 1 NR2 $T=424700 719160 1 0 $X=424700 $Y=713740
X3744 2196 2 2377 2342 1 NR2 $T=425320 678840 1 0 $X=425320 $Y=673420
X3745 2259 2 2378 236 1 NR2 $T=429660 668760 0 180 $X=427800 $Y=663340
X3746 2383 2 2379 2317 1 NR2 $T=429660 678840 1 180 $X=427800 $Y=678460
X3747 2254 2 2374 222 1 NR2 $T=429660 719160 0 180 $X=427800 $Y=713740
X3748 2372 2 2393 2352 1 NR2 $T=430280 557880 1 180 $X=428420 $Y=557500
X3749 2259 2 2384 222 1 NR2 $T=430280 678840 0 180 $X=428420 $Y=673420
X3750 2254 2 2382 2342 1 NR2 $T=429040 699000 1 0 $X=429040 $Y=693580
X3751 2316 2 2400 2333 1 NR2 $T=430900 578040 1 0 $X=430900 $Y=572620
X3752 198 2 250 249 1 NR2 $T=435860 719160 0 0 $X=435860 $Y=718780
X3753 198 2 2437 233 1 NR2 $T=440820 709080 0 180 $X=438960 $Y=703660
X3754 2368 2 251 2433 1 NR2 $T=441440 547800 0 180 $X=439580 $Y=542380
X3755 2143 2 2434 233 1 NR2 $T=441440 688920 1 180 $X=439580 $Y=688540
X3756 2436 2 2463 2366 1 NR2 $T=444540 658680 1 180 $X=442680 $Y=658300
X3757 2383 2 2471 2227 1 NR2 $T=442680 688920 0 0 $X=442680 $Y=688540
X3758 2436 2 2480 2227 1 NR2 $T=443300 668760 1 0 $X=443300 $Y=663340
X3759 2383 2 2452 2366 1 NR2 $T=445160 668760 1 180 $X=443300 $Y=668380
X3760 254 2 2477 256 1 NR2 $T=443300 678840 0 0 $X=443300 $Y=678460
X3761 2143 2 2488 249 1 NR2 $T=443300 688920 1 0 $X=443300 $Y=683500
X3762 2420 2 2476 2227 1 NR2 $T=446400 658680 1 180 $X=444540 $Y=658300
X3763 254 2 2511 2544 1 NR2 $T=449500 678840 1 0 $X=449500 $Y=673420
X3764 224 2 265 245 1 NR2 $T=451980 719160 0 0 $X=451980 $Y=718780
X3765 2514 2 2533 256 1 NR2 $T=455080 699000 0 180 $X=453220 $Y=693580
X3766 2528 2 2529 256 1 NR2 $T=455080 709080 1 180 $X=453220 $Y=708700
X3767 2436 2 2523 268 1 NR2 $T=453840 547800 0 0 $X=453840 $Y=547420
X3768 279 2 2522 2485 1 NR2 $T=455700 699000 1 180 $X=453840 $Y=698620
X3769 2460 2 2551 245 1 NR2 $T=455700 688920 1 0 $X=455700 $Y=683500
X3770 2514 2 2552 253 1 NR2 $T=455700 699000 1 0 $X=455700 $Y=693580
X3771 268 2 2537 2420 1 NR2 $T=456940 547800 0 0 $X=456940 $Y=547420
X3772 2460 2 2554 253 1 NR2 $T=458800 658680 0 180 $X=456940 $Y=653260
X3773 183 2 2534 2544 1 NR2 $T=456940 719160 0 0 $X=456940 $Y=718780
X3774 2143 2 2549 245 1 NR2 $T=459420 668760 1 180 $X=457560 $Y=668380
X3775 2528 2 2550 2516 1 NR2 $T=457560 678840 0 0 $X=457560 $Y=678460
X3776 2266 2 2568 2391 1 NR2 $T=461280 658680 0 180 $X=459420 $Y=653260
X3777 281 2 274 2544 1 NR2 $T=463760 719160 1 180 $X=461900 $Y=718780
X3778 276 2 2525 2588 1 NR2 $T=462520 547800 0 0 $X=462520 $Y=547420
X3779 2577 2 2566 277 1 NR2 $T=462520 578040 0 0 $X=462520 $Y=577660
X3780 2266 2 2585 2414 1 NR2 $T=462520 648600 1 0 $X=462520 $Y=643180
X3781 2565 2 2582 2588 1 NR2 $T=463140 557880 0 0 $X=463140 $Y=557500
X3782 2584 2 2594 282 1 NR2 $T=463760 567960 0 0 $X=463760 $Y=567580
X3783 2584 2 2592 268 1 NR2 $T=464380 547800 1 0 $X=464380 $Y=542380
X3784 2383 2 2567 277 1 NR2 $T=466240 578040 1 180 $X=464380 $Y=577660
X3785 2593 2 2616 2565 1 NR2 $T=465620 567960 1 0 $X=465620 $Y=562540
X3786 2577 2 2580 282 1 NR2 $T=467480 578040 0 180 $X=465620 $Y=572620
X3787 280 2 2596 2588 1 NR2 $T=466240 547800 0 0 $X=466240 $Y=547420
X3788 2612 2 2610 2346 1 NR2 $T=468100 638520 0 180 $X=466240 $Y=633100
X3789 2611 2 2603 2414 1 NR2 $T=468100 648600 0 180 $X=466240 $Y=643180
X3790 2611 2 2598 2346 1 NR2 $T=468100 648600 1 180 $X=466240 $Y=648220
X3791 279 2 2629 2516 1 NR2 $T=466240 699000 0 0 $X=466240 $Y=698620
X3792 280 2 2570 2593 1 NR2 $T=466860 547800 1 0 $X=466860 $Y=542380
X3793 276 2 2595 2593 1 NR2 $T=466860 557880 1 0 $X=466860 $Y=552460
X3794 2383 2 2562 2613 1 NR2 $T=467480 578040 0 0 $X=467480 $Y=577660
X3795 2617 2 2608 2565 1 NR2 $T=469960 557880 1 180 $X=468100 $Y=557500
X3796 2630 2 2563 2617 1 NR2 $T=471820 557880 0 180 $X=469960 $Y=552460
X3797 2460 2 2649 2588 1 NR2 $T=471200 598200 1 0 $X=471200 $Y=592780
X3798 2577 2 2631 2588 1 NR2 $T=473680 578040 0 180 $X=471820 $Y=572620
X3799 280 2 2639 2617 1 NR2 $T=473060 557880 1 0 $X=473060 $Y=552460
X3800 2630 2 2632 2593 1 NR2 $T=473680 547800 0 0 $X=473680 $Y=547420
X3801 276 2 2638 282 1 NR2 $T=474920 547800 1 0 $X=474920 $Y=542380
X3802 2658 2 2667 282 1 NR2 $T=480500 567960 0 180 $X=478640 $Y=562540
X3803 2584 2 2674 2593 1 NR2 $T=480500 547800 0 0 $X=480500 $Y=547420
X3804 2584 2 2675 2588 1 NR2 $T=482360 557880 0 180 $X=480500 $Y=552460
X3805 2630 2 2643 306 1 NR2 $T=481120 557880 0 0 $X=481120 $Y=557500
X3806 2617 2 2682 2671 1 NR2 $T=482360 557880 1 0 $X=482360 $Y=552460
X3807 2678 2 2679 2617 1 NR2 $T=482360 567960 1 0 $X=482360 $Y=562540
X3808 306 2 2695 2565 1 NR2 $T=486080 557880 1 180 $X=484220 $Y=557500
X3809 2593 2 2706 2671 1 NR2 $T=485460 557880 1 0 $X=485460 $Y=552460
X3810 2698 2 2702 317 1 NR2 $T=485460 567960 1 0 $X=485460 $Y=562540
X3811 2528 2 2699 306 1 NR2 $T=487320 567960 1 180 $X=485460 $Y=567580
X3812 2436 2 2700 2613 1 NR2 $T=489180 588120 0 180 $X=487320 $Y=582700
X3813 2528 2 2718 317 1 NR2 $T=488560 557880 0 0 $X=488560 $Y=557500
X3814 306 2 2748 2671 1 NR2 $T=492900 557880 0 180 $X=491040 $Y=552460
X3815 2565 2 2732 321 1 NR2 $T=491040 557880 0 0 $X=491040 $Y=557500
X3816 2725 2 2733 2266 1 NR2 $T=491040 578040 1 0 $X=491040 $Y=572620
X3817 2725 2 2769 2420 1 NR2 $T=496620 578040 0 180 $X=494760 $Y=572620
X3818 2678 2 2772 321 1 NR2 $T=497860 567960 0 180 $X=496000 $Y=562540
X3819 2782 2 2755 2633 1 NR2 $T=497860 567960 1 180 $X=496000 $Y=567580
X3820 2613 2 2765 2619 1 NR2 $T=496000 588120 0 0 $X=496000 $Y=587740
X3821 306 2 2791 2658 1 NR2 $T=497860 567960 1 0 $X=497860 $Y=562540
X3822 2617 2 2792 2764 1 NR2 $T=498480 557880 0 0 $X=498480 $Y=557500
X3823 2782 2 330 2611 1 NR2 $T=499720 547800 1 0 $X=499720 $Y=542380
X3824 2802 2 2799 2658 1 NR2 $T=503440 557880 1 180 $X=501580 $Y=557500
X3825 2420 2 2815 298 1 NR2 $T=504680 578040 1 0 $X=504680 $Y=572620
X3826 2834 2 2835 321 1 NR2 $T=508400 547800 0 180 $X=506540 $Y=542380
X3827 317 2 2829 2658 1 NR2 $T=507160 557880 1 0 $X=507160 $Y=552460
X3828 2727 2 2836 2802 1 NR2 $T=509020 567960 0 180 $X=507160 $Y=562540
X3829 2727 2 2837 298 1 NR2 $T=509020 578040 0 180 $X=507160 $Y=572620
X3830 2613 2 2841 2266 1 NR2 $T=507160 588120 0 0 $X=507160 $Y=587740
X3831 2834 2 349 350 1 NR2 $T=508400 547800 1 0 $X=508400 $Y=542380
X3832 2789 2 2843 2658 1 NR2 $T=510260 547800 1 180 $X=508400 $Y=547420
X3833 344 2 2846 350 1 NR2 $T=509020 537720 0 0 $X=509020 $Y=537340
X3834 2633 2 2850 300 1 NR2 $T=509020 578040 1 0 $X=509020 $Y=572620
X3835 2678 2 2847 350 1 NR2 $T=509640 557880 0 0 $X=509640 $Y=557500
X3836 344 2 356 2876 1 NR2 $T=513980 537720 0 0 $X=513980 $Y=537340
X3837 2420 2 2854 300 1 NR2 $T=513980 578040 1 0 $X=513980 $Y=572620
X3838 2633 2 2872 360 1 NR2 $T=513980 578040 0 0 $X=513980 $Y=577660
X3839 2725 2 2890 2611 1 NR2 $T=517700 547800 0 180 $X=515840 $Y=542380
X3840 2619 2 2879 360 1 NR2 $T=517700 588120 0 180 $X=515840 $Y=582700
X3841 2834 2 2893 2876 1 NR2 $T=519560 537720 1 180 $X=517700 $Y=537340
X3842 2782 2 2880 2612 1 NR2 $T=518940 557880 0 0 $X=518940 $Y=557500
X3843 2727 2 2910 300 1 NR2 $T=520800 578040 1 0 $X=520800 $Y=572620
X3844 2782 2 2903 2920 1 NR2 $T=521420 557880 0 0 $X=521420 $Y=557500
X3845 2725 2 2926 2619 1 NR2 $T=521420 567960 0 0 $X=521420 $Y=567580
X3846 2613 2 2921 2633 1 NR2 $T=521420 588120 1 0 $X=521420 $Y=582700
X3847 2725 2 2938 2633 1 NR2 $T=523280 578040 1 0 $X=523280 $Y=572620
X3848 2782 2 2943 2619 1 NR2 $T=526380 557880 0 0 $X=526380 $Y=557500
X3849 2727 2 2952 360 1 NR2 $T=528240 578040 0 180 $X=526380 $Y=572620
X3850 425 2 3152 3155 1 NR2 $T=567300 547800 1 0 $X=567300 $Y=542380
X3851 471 2 3179 3182 1 NR2 $T=574740 557880 1 180 $X=572880 $Y=557500
X3852 3070 2 3139 3192 1 NR2 $T=572880 567960 0 0 $X=572880 $Y=567580
X3853 462 2 3191 3192 1 NR2 $T=572880 578040 1 0 $X=572880 $Y=572620
X3854 3148 2 3193 474 1 NR2 $T=573500 567960 1 0 $X=573500 $Y=562540
X3855 471 2 3196 3155 1 NR2 $T=575980 537720 1 180 $X=574120 $Y=537340
X3856 426 2 3202 413 1 NR2 $T=574120 547800 0 0 $X=574120 $Y=547420
X3857 3155 2 3199 3070 1 NR2 $T=576600 578040 0 180 $X=574740 $Y=572620
X3858 3203 2 3198 2920 1 NR2 $T=576600 557880 0 0 $X=576600 $Y=557500
X3859 471 2 483 2920 1 NR2 $T=579080 557880 0 0 $X=579080 $Y=557500
X3860 471 2 3232 413 1 NR2 $T=583420 557880 1 180 $X=581560 $Y=557500
X3861 3070 2 3247 3220 1 NR2 $T=587140 578040 1 0 $X=587140 $Y=572620
X3862 426 2 3244 512 1 NR2 $T=588380 557880 1 0 $X=588380 $Y=552460
X3863 3203 2 3267 3182 1 NR2 $T=588380 567960 1 0 $X=588380 $Y=562540
X3864 497 2 3271 512 1 NR2 $T=589000 547800 1 0 $X=589000 $Y=542380
X3865 3070 2 3276 3182 1 NR2 $T=590240 578040 1 0 $X=590240 $Y=572620
X3866 3024 2 3324 3182 1 NR2 $T=601400 567960 1 180 $X=599540 $Y=567580
X3867 3024 2 3297 3155 1 NR2 $T=599540 578040 1 0 $X=599540 $Y=572620
X3868 3321 2 3328 512 1 NR2 $T=600780 547800 0 0 $X=600780 $Y=547420
X3869 3330 2 3332 3148 1 NR2 $T=602640 588120 1 0 $X=602640 $Y=582700
X3870 3024 2 3347 3350 1 NR2 $T=605120 578040 1 0 $X=605120 $Y=572620
X3871 552 2 3376 3363 1 NR2 $T=607600 547800 0 0 $X=607600 $Y=547420
X3872 3203 2 3371 3363 1 NR2 $T=608220 567960 1 0 $X=608220 $Y=562540
X3873 3203 2 3362 3350 1 NR2 $T=608220 567960 0 0 $X=608220 $Y=567580
X3874 406 2 3381 559 1 NR2 $T=608840 537720 0 0 $X=608840 $Y=537340
X3875 3364 2 3382 537 1 NR2 $T=610080 588120 1 0 $X=610080 $Y=582700
X3876 3364 2 3403 3220 1 NR2 $T=615040 578040 0 180 $X=613180 $Y=572620
X3877 537 2 3392 474 1 NR2 $T=615660 567960 0 180 $X=613800 $Y=562540
X3878 565 2 3411 474 1 NR2 $T=615040 547800 0 0 $X=615040 $Y=547420
X3879 537 2 3415 3148 1 NR2 $T=616900 578040 1 0 $X=616900 $Y=572620
X3880 3396 2 2924 3454 1 NR2 $T=622480 658680 0 0 $X=622480 $Y=658300
X3881 593 2 3396 3429 1 NR2 $T=624340 678840 0 180 $X=622480 $Y=673420
X3882 3434 2 3442 3421 1 NR2 $T=626200 699000 0 180 $X=624340 $Y=693580
X3883 3459 2 3460 3450 1 NR2 $T=626820 588120 1 180 $X=624960 $Y=587740
X3884 3457 2 3454 3468 1 NR2 $T=626200 658680 0 0 $X=626200 $Y=658300
X3885 3434 2 3498 3505 1 NR2 $T=632400 688920 1 0 $X=632400 $Y=683500
X3886 2669 2 3513 3432 1 NR2 $T=633020 709080 1 0 $X=633020 $Y=703660
X3887 3485 2 3532 3497 1 NR2 $T=636740 578040 0 0 $X=636740 $Y=577660
X3888 3527 2 3610 3579 1 NR2 $T=651000 709080 0 180 $X=649140 $Y=703660
X3889 668 2 3452 3726 1 NR2 $T=674560 699000 1 180 $X=672700 $Y=698620
X3890 718 2 3954 3503 1 NR2 $T=717960 709080 1 180 $X=716100 $Y=708700
X3891 3954 2 720 3706 1 NR2 $T=718580 719160 1 0 $X=718580 $Y=713740
X3892 3995 2 3984 3005 1 NR2 $T=724780 719160 1 0 $X=724780 $Y=713740
X3893 3005 2 4006 3998 1 NR2 $T=727260 719160 1 180 $X=725400 $Y=718780
X3894 4006 2 4008 727 1 NR2 $T=727260 719160 0 0 $X=727260 $Y=718780
X3895 733 2 4022 4024 1 NR2 $T=733460 578040 1 180 $X=731600 $Y=577660
X3896 4027 2 4034 739 1 NR2 $T=732840 648600 0 0 $X=732840 $Y=648220
X3897 4027 2 4029 4024 1 NR2 $T=733460 628440 0 0 $X=733460 $Y=628060
X3898 735 2 4030 4024 1 NR2 $T=735320 648600 0 180 $X=733460 $Y=643180
X3899 734 2 4021 4049 1 NR2 $T=734700 719160 1 0 $X=734700 $Y=713740
X3900 4046 2 4050 743 1 NR2 $T=735940 588120 0 0 $X=735940 $Y=587740
X3901 745 2 4051 4024 1 NR2 $T=737800 608280 1 180 $X=735940 $Y=607900
X3902 4046 2 3985 4024 1 NR2 $T=738420 598200 0 180 $X=736560 $Y=592780
X3903 744 2 4053 4060 1 NR2 $T=737180 608280 1 0 $X=737180 $Y=602860
X3904 746 2 750 743 1 NR2 $T=737800 537720 0 0 $X=737800 $Y=537340
X3905 744 2 4039 4046 1 NR2 $T=739660 618360 0 180 $X=737800 $Y=612940
X3906 757 2 4055 4049 1 NR2 $T=741520 709080 0 180 $X=739660 $Y=703660
X3907 754 2 4052 4049 1 NR2 $T=739660 709080 0 0 $X=739660 $Y=708700
X3908 4060 2 4069 743 1 NR2 $T=743380 588120 0 180 $X=741520 $Y=582700
X3909 4077 2 4072 760 1 NR2 $T=741520 688920 0 0 $X=741520 $Y=688540
X3910 4027 2 4083 760 1 NR2 $T=744620 688920 0 180 $X=742760 $Y=683500
X3911 761 2 4091 763 1 NR2 $T=742760 709080 0 0 $X=742760 $Y=708700
X3912 775 2 4156 763 1 NR2 $T=755780 709080 0 0 $X=755780 $Y=708700
X3913 778 2 4168 4157 1 NR2 $T=758260 638520 1 180 $X=756400 $Y=638140
X3914 4164 2 4080 4157 1 NR2 $T=757020 668760 1 0 $X=757020 $Y=663340
X3915 4164 2 4176 779 1 NR2 $T=757640 688920 1 0 $X=757640 $Y=683500
X3916 4184 2 3978 763 1 NR2 $T=761360 668760 1 180 $X=759500 $Y=668380
X3917 4184 2 4180 779 1 NR2 $T=762600 678840 1 180 $X=760740 $Y=678460
X3918 786 2 4148 4157 1 NR2 $T=764460 638520 1 180 $X=762600 $Y=638140
X3919 784 2 4110 789 1 NR2 $T=762600 719160 0 0 $X=762600 $Y=718780
X3920 4223 2 794 782 1 NR2 $T=771280 719160 0 0 $X=771280 $Y=718780
X3921 788 2 806 805 1 NR2 $T=781820 719160 1 180 $X=779960 $Y=718780
X3922 4027 2 4540 858 1 NR2 $T=825220 688920 0 0 $X=825220 $Y=688540
X3923 4077 2 4522 858 1 NR2 $T=828320 709080 0 180 $X=826460 $Y=703660
X3924 4184 2 4534 867 1 NR2 $T=832660 699000 1 0 $X=832660 $Y=693580
X3925 4060 2 4564 862 1 NR2 $T=835140 588120 0 0 $X=835140 $Y=587740
X3926 4046 2 4585 862 1 NR2 $T=837620 598200 1 180 $X=835760 $Y=597820
X3927 4164 2 4523 867 1 NR2 $T=838240 699000 1 0 $X=838240 $Y=693580
X3928 4184 2 4566 876 1 NR2 $T=839480 668760 1 0 $X=839480 $Y=663340
X3929 4164 2 4561 876 1 NR2 $T=839480 678840 1 0 $X=839480 $Y=673420
X3930 4027 2 4615 878 1 NR2 $T=840100 688920 1 0 $X=840100 $Y=683500
X3931 880 2 4588 4164 1 NR2 $T=842580 658680 1 180 $X=840720 $Y=658300
X3932 4164 2 4630 843 1 NR2 $T=842580 658680 0 0 $X=842580 $Y=658300
X3933 4077 2 4685 803 1 NR2 $T=854360 658680 0 0 $X=854360 $Y=658300
X3934 4060 2 4742 890 1 NR2 $T=862420 598200 0 180 $X=860560 $Y=592780
X3935 4652 2 4751 890 1 NR2 $T=864900 598200 0 180 $X=863040 $Y=592780
X3936 735 2 4809 810 1 NR2 $T=872960 658680 1 0 $X=872960 $Y=653260
X3937 4617 2 4852 810 1 NR2 $T=881640 628440 0 180 $X=879780 $Y=623020
X3938 733 2 4848 928 1 NR2 $T=883500 588120 0 180 $X=881640 $Y=582700
X3939 4652 2 4898 928 1 NR2 $T=889080 588120 0 180 $X=887220 $Y=582700
X3940 4060 2 5369 1020 1 NR2 $T=971540 588120 1 0 $X=971540 $Y=582700
X3941 4617 2 5360 1031 1 NR2 $T=974020 688920 0 0 $X=974020 $Y=688540
X3942 4617 2 5372 803 1 NR2 $T=978980 628440 0 180 $X=977120 $Y=623020
X3943 4652 2 5393 1020 1 NR2 $T=982080 588120 0 180 $X=980220 $Y=582700
X3944 880 2 5402 1038 1 NR2 $T=982080 668760 1 0 $X=982080 $Y=663340
X3945 735 2 5441 1045 1 NR2 $T=985180 678840 0 0 $X=985180 $Y=678460
X3946 4617 2 5453 1045 1 NR2 $T=986420 658680 1 0 $X=986420 $Y=653260
X3947 4652 2 5457 1061 1 NR2 $T=988280 588120 1 0 $X=988280 $Y=582700
X3948 733 2 5470 1061 1 NR2 $T=993860 588120 0 180 $X=992000 $Y=582700
X3949 1038 2 5482 876 1 NR2 $T=993860 668760 0 0 $X=993860 $Y=668380
X3950 876 2 5483 1053 1 NR2 $T=996960 668760 0 0 $X=996960 $Y=668380
X3951 1048 2 5534 1053 1 NR2 $T=996960 688920 0 0 $X=996960 $Y=688540
X3952 4652 2 5521 1068 1 NR2 $T=1000680 598200 0 180 $X=998820 $Y=592780
X3953 1960 12 1 2 INV12CK $T=354020 628440 0 180 $X=344100 $Y=623020
X3954 1960 136 1 2 INV12CK $T=398660 618360 0 0 $X=398660 $Y=617980
X3955 700 3860 1 2 INV12CK $T=698740 638520 0 0 $X=698740 $Y=638140
X3956 4047 3292 1 2 INV12CK $T=736560 598200 0 180 $X=726640 $Y=592780
X3957 4047 553 1 2 INV12CK $T=740280 578040 0 0 $X=740280 $Y=577660
X3958 815 4047 1 2 INV12CK $T=797940 578040 0 0 $X=797940 $Y=577660
X3959 4047 839 1 2 INV12CK $T=812820 588120 0 0 $X=812820 $Y=587740
X3960 4281 4570 1 2 INV12CK $T=829560 709080 0 0 $X=829560 $Y=708700
X3961 4570 837 1 2 INV12CK $T=877300 719160 0 180 $X=867380 $Y=713740
X3962 3860 982 1 2 INV12CK $T=922560 547800 0 0 $X=922560 $Y=547420
X3963 4570 970 1 2 INV12CK $T=938680 719160 0 180 $X=928760 $Y=713740
X3964 5370 969 1 2 INV12CK $T=977740 547800 0 180 $X=967820 $Y=542380
X3965 5370 4818 1 2 INV12CK $T=983320 567960 0 180 $X=973400 $Y=562540
X3966 5370 1025 1 2 INV12CK $T=992000 557880 0 0 $X=992000 $Y=557500
X3967 4570 1098 1 2 INV12CK $T=1012460 719160 0 0 $X=1012460 $Y=718780
X3968 1157 1121 1 2 INV12CK $T=1085620 557880 0 180 $X=1075700 $Y=552460
X3969 1157 5560 1 2 INV12CK $T=1085620 578040 0 180 $X=1075700 $Y=572620
X3970 5425 1157 1 2 INV12CK $T=1078800 547800 1 0 $X=1078800 $Y=542380
X3971 33 32 2 1 35 OR2 $T=241800 719160 1 0 $X=241800 $Y=713740
X3972 1690 1684 2 1 1677 OR2 $T=301940 547800 1 180 $X=299460 $Y=547420
X3973 98 122 2 1 114 OR2 $T=313720 537720 1 180 $X=311240 $Y=537340
X3974 1971 1841 2 1 1948 OR2 $T=355880 678840 0 0 $X=355880 $Y=678460
X3975 2290 2321 2 1 2332 OR2 $T=419740 547800 0 0 $X=419740 $Y=547420
X3976 2331 2287 2 1 2355 OR2 $T=423460 578040 1 0 $X=423460 $Y=572620
X3977 2327 2300 2 1 2361 OR2 $T=429040 557880 0 180 $X=426560 $Y=552460
X3978 2411 2286 2 1 2427 OR2 $T=435860 557880 1 0 $X=435860 $Y=552460
X3979 292 299 2 1 260 OR2 $T=480500 719160 1 180 $X=478020 $Y=718780
X3980 458 497 2 1 3252 OR2 $T=589000 547800 0 180 $X=586520 $Y=542380
X3981 3295 3269 2 1 3237 OR2 $T=592720 648600 1 180 $X=590240 $Y=648220
X3982 3296 3297 2 1 3300 OR2 $T=598920 578040 1 180 $X=596440 $Y=577660
X3983 458 426 2 1 3335 OR2 $T=601400 547800 1 0 $X=601400 $Y=542380
X3984 458 3321 2 1 3352 OR2 $T=605120 547800 0 0 $X=605120 $Y=547420
X3985 458 3203 2 1 3375 OR2 $T=606360 547800 1 0 $X=606360 $Y=542380
X3986 3480 3434 2 1 3466 OR2 $T=630540 688920 0 180 $X=628060 $Y=683500
X3987 3516 619 2 1 3546 OR2 $T=636120 588120 1 0 $X=636120 $Y=582700
X3988 3511 619 2 1 3464 OR2 $T=636120 598200 1 0 $X=636120 $Y=592780
X3989 739 4077 2 1 3824 OR2 $T=743380 678840 0 180 $X=740900 $Y=673420
X3990 4129 777 2 1 782 OR2 $T=758880 719160 0 0 $X=758880 $Y=718780
X3991 789 788 2 1 4049 OR2 $T=765080 719160 0 180 $X=762600 $Y=713740
X3992 792 784 2 1 803 OR2 $T=776860 719160 0 0 $X=776860 $Y=718780
X3993 792 788 2 1 810 OR2 $T=781820 719160 0 0 $X=781820 $Y=718780
X3994 881 4060 2 1 4609 OR2 $T=843200 598200 1 180 $X=840720 $Y=597820
X3995 881 4046 2 1 869 OR2 $T=843820 588120 0 0 $X=843820 $Y=587740
X3996 884 4617 2 1 4562 OR2 $T=846920 648600 1 180 $X=844440 $Y=648220
X3997 884 4077 2 1 4672 OR2 $T=849400 658680 0 0 $X=849400 $Y=658300
X3998 878 4077 2 1 4673 OR2 $T=849400 668760 1 0 $X=849400 $Y=663340
X3999 1036 735 2 1 5379 OR2 $T=981460 678840 0 0 $X=981460 $Y=678460
X4000 1031 735 2 1 5442 OR2 $T=984560 709080 0 0 $X=984560 $Y=708700
X4001 1036 4617 2 1 5385 OR2 $T=986420 658680 0 0 $X=986420 $Y=658300
X4002 1036 1073 2 1 1075 OR2 $T=994480 719160 0 0 $X=994480 $Y=718780
X4003 1076 733 2 1 5494 OR2 $T=996960 598200 0 0 $X=996960 $Y=597820
X4004 1511 1518 1 2 1520 AN2 $T=274040 547800 1 180 $X=271560 $Y=547420
X4005 1743 1744 1 2 1757 AN2 $T=311860 567960 1 0 $X=311860 $Y=562540
X4006 1886 1877 1 2 1870 AN2 $T=340380 567960 1 180 $X=337900 $Y=567580
X4007 1995 1977 1 2 1986 AN2 $T=363320 578040 1 180 $X=360840 $Y=577660
X4008 2014 1945 1 2 1985 AN2 $T=368900 618360 1 180 $X=366420 $Y=617980
X4009 2228 218 1 2 219 AN2 $T=406720 547800 1 0 $X=406720 $Y=542380
X4010 2206 218 1 2 2261 AN2 $T=409200 547800 1 0 $X=409200 $Y=542380
X4011 2220 2256 1 2 2263 AN2 $T=409200 557880 0 0 $X=409200 $Y=557500
X4012 2242 2256 1 2 2278 AN2 $T=409200 567960 0 0 $X=409200 $Y=567580
X4013 2247 2256 1 2 2302 AN2 $T=416640 557880 1 0 $X=416640 $Y=552460
X4014 375 368 1 2 2929 AN2 $T=527000 537720 1 180 $X=524520 $Y=537340
X4015 3275 506 1 2 3283 AN2 $T=590240 709080 1 0 $X=590240 $Y=703660
X4016 3285 508 1 2 3212 AN2 $T=592720 719160 0 180 $X=590240 $Y=713740
X4017 3285 516 1 2 3189 AN2 $T=595820 719160 0 180 $X=593340 $Y=713740
X4018 3285 517 1 2 3229 AN2 $T=596440 709080 0 180 $X=593960 $Y=703660
X4019 3275 518 1 2 3269 AN2 $T=596440 709080 1 180 $X=593960 $Y=708700
X4020 3285 521 1 2 3250 AN2 $T=598300 719160 0 180 $X=595820 $Y=713740
X4021 3285 531 1 2 3261 AN2 $T=601400 719160 0 180 $X=598920 $Y=713740
X4022 3285 535 1 2 3306 AN2 $T=600780 709080 0 0 $X=600780 $Y=708700
X4023 3429 3395 1 2 3436 AN2 $T=620000 678840 1 0 $X=620000 $Y=673420
X4024 3275 595 1 2 3412 AN2 $T=625580 709080 0 180 $X=623100 $Y=703660
X4025 3275 597 1 2 3444 AN2 $T=626200 699000 1 180 $X=623720 $Y=698620
X4026 3275 598 1 2 3438 AN2 $T=628680 709080 0 180 $X=626200 $Y=703660
X4027 3541 627 1 2 3531 AN2 $T=642320 699000 1 180 $X=639840 $Y=698620
X4028 17 2 1244 16 1266 1 NR3 $T=225060 719160 1 180 $X=221960 $Y=718780
X4029 1310 2 28 1340 1305 1 NR3 $T=234980 719160 0 0 $X=234980 $Y=718780
X4030 1324 2 32 1333 1291 1 NR3 $T=240560 699000 0 0 $X=240560 $Y=698620
X4031 1612 1705 1 1801 2 OR2B1S $T=319920 567960 1 0 $X=319920 $Y=562540
X4032 1612 1816 1 1836 2 OR2B1S $T=332320 557880 0 180 $X=329220 $Y=552460
X4033 2039 2071 1 2150 2 OR2B1S $T=388740 557880 0 0 $X=388740 $Y=557500
X4034 2039 2065 1 2232 2 OR2B1S $T=401760 578040 1 0 $X=401760 $Y=572620
X4035 2573 2641 1 2672 2 OR2B1S $T=478020 618360 0 0 $X=478020 $Y=617980
X4036 2807 2787 1 2745 2 OR2B1S $T=505920 658680 1 180 $X=502820 $Y=658300
X4037 2807 3031 1 3037 2 OR2B1S $T=546220 668760 0 180 $X=543120 $Y=663340
X4038 3032 3038 1 3052 2 OR2B1S $T=544360 567960 0 0 $X=544360 $Y=567580
X4039 3032 3096 1 3130 2 OR2B1S $T=559240 547800 0 0 $X=559240 $Y=547420
X4040 3188 3156 1 3153 2 OR2B1S $T=574120 648600 0 180 $X=571020 $Y=643180
X4041 3219 3151 1 3230 2 OR2B1S $T=582800 608280 1 0 $X=582800 $Y=602860
X4042 3188 3207 1 3268 2 OR2B1S $T=591480 618360 1 0 $X=591480 $Y=612940
X4043 592 3369 1 3428 2 OR2B1S $T=624340 598200 0 180 $X=621240 $Y=592780
X4044 3432 2669 1 587 2 OR2B1S $T=632400 709080 0 180 $X=629300 $Y=703660
X4045 3533 3527 1 3421 2 OR2B1S $T=638600 699000 0 180 $X=635500 $Y=693580
X4046 5358 5499 1 5516 2 OR2B1S $T=997580 648600 0 0 $X=997580 $Y=648220
X4047 2886 1 2 2915 396 311 384 382 1233 ICV_8 $T=523280 719160 0 0 $X=523280 $Y=718780
X4048 2937 1 2 3012 3013 385 393 3019 1233 ICV_8 $T=535060 557880 1 0 $X=535060 $Y=552460
X4049 404 1 2 411 3105 311 3017 3059 1233 ICV_8 $T=543120 688920 0 0 $X=543120 $Y=688540
X4050 3821 1 2 3846 3893 3292 3750 3850 1233 ICV_8 $T=689440 608280 0 0 $X=689440 $Y=607900
X4051 3917 1 2 3943 3971 724 3912 3917 1233 ICV_8 $T=710520 658680 1 0 $X=710520 $Y=653260
X4052 3930 1 2 3957 4012 553 3876 633 1233 ICV_8 $T=713000 547800 1 0 $X=713000 $Y=542380
X4053 4162 1 2 4138 4243 724 4133 3483 1233 ICV_8 $T=758260 648600 0 0 $X=758260 $Y=648220
X4054 4264 1 2 4289 4331 742 4278 4264 1233 ICV_8 $T=776860 598200 1 0 $X=776860 $Y=592780
X4055 4367 1 2 4386 4413 724 4217 3435 1233 ICV_8 $T=797320 668760 1 0 $X=797320 $Y=663340
X4056 4382 1 2 4397 4384 724 4417 3462 1233 ICV_8 $T=800420 638520 1 0 $X=800420 $Y=633100
X4057 4399 1 2 4414 4429 837 4390 4399 1233 ICV_8 $T=802280 699000 1 0 $X=802280 $Y=693580
X4058 4371 1 2 4422 4436 839 4420 4371 1233 ICV_8 $T=802900 567960 1 0 $X=802900 $Y=562540
X4059 921 1 2 926 4907 837 4805 4846 1233 ICV_8 $T=875440 709080 1 0 $X=875440 $Y=703660
X4060 5018 1 2 5056 5088 970 4902 5010 1233 ICV_8 $T=910780 658680 1 0 $X=910780 $Y=653260
X4061 5098 1 2 5129 5197 970 5127 5134 1233 ICV_8 $T=924420 709080 0 0 $X=924420 $Y=708700
X4062 5163 1 2 5156 5294 970 5243 5254 1233 ICV_8 $T=944260 658680 1 0 $X=944260 $Y=653260
X4063 5232 1 2 5256 5286 970 5255 5237 1233 ICV_8 $T=946120 678840 0 0 $X=946120 $Y=678460
X4064 5244 1 2 5272 5305 4818 5243 5244 1233 ICV_8 $T=947360 628440 0 0 $X=947360 $Y=628060
X4065 5192 1 2 5234 5378 1025 5288 5336 1233 ICV_8 $T=963480 557880 0 0 $X=963480 $Y=557500
X4066 5636 1 2 5664 5718 5560 5683 5667 1233 ICV_8 $T=1019900 628440 1 0 $X=1019900 $Y=623020
X4067 5847 1 2 5851 5919 5560 5683 5871 1233 ICV_8 $T=1057720 608280 1 0 $X=1057720 $Y=602860
X4068 5953 1 2 5963 6033 5560 5962 5974 1233 ICV_8 $T=1078800 618360 0 0 $X=1078800 $Y=617980
X4069 1169 1 2 6078 6124 1098 5936 1169 1233 ICV_8 $T=1097400 719160 1 0 $X=1097400 $Y=713740
X4070 1181 1 2 6134 6141 1098 1175 6098 1233 ICV_8 $T=1107940 709080 0 0 $X=1107940 $Y=708700
X4071 6128 1 2 6115 6180 1098 6178 6129 1233 ICV_8 $T=1112280 658680 0 0 $X=1112280 $Y=658300
X4072 3875 3713 2 1 3894 3458 3771 3760 3854 3864 3779 1233 ICV_9 $T=695020 688920 1 0 $X=695020 $Y=683500
X4073 4135 4075 2 1 4171 785 4134 774 4172 4114 3710 1233 ICV_9 $T=757640 567960 0 0 $X=757640 $Y=567580
X4074 4345 4079 2 1 4366 4357 4025 4106 4297 4339 3484 1233 ICV_9 $T=788640 608280 0 0 $X=788640 $Y=607900
X4075 3517 4041 2 1 4418 4357 4025 4106 4372 4381 3380 1233 ICV_9 $T=797320 608280 0 0 $X=797320 $Y=607900
X4076 4863 4822 2 1 4932 816 4795 4884 4640 4894 4832 1233 ICV_9 $T=887220 638520 0 0 $X=887220 $Y=638140
X4077 5036 4880 2 1 5059 4950 4690 4703 4972 5012 5017 1233 ICV_9 $T=908300 688920 1 0 $X=908300 $Y=683500
X4078 5216 5207 2 1 5242 5155 5170 5021 5054 5203 5187 1233 ICV_9 $T=939920 618360 1 0 $X=939920 $Y=612940
X4079 5272 4955 2 1 5305 5280 5091 5159 5230 5244 5263 1233 ICV_9 $T=948600 638520 1 0 $X=948600 $Y=633100
X4080 5601 5494 2 1 5624 5445 5543 5496 5524 5570 5555 1233 ICV_9 $T=1009980 608280 1 0 $X=1009980 $Y=602860
X4081 5784 5579 2 1 5790 5797 5681 5460 5739 5756 5757 1233 ICV_9 $T=1042840 668760 1 0 $X=1042840 $Y=663340
X4082 5791 5794 2 1 5820 1097 5502 5777 5730 1124 5768 1233 ICV_9 $T=1044700 547800 0 0 $X=1044700 $Y=547420
X4083 5893 5826 2 1 5916 5910 5680 5745 5855 5871 5886 1233 ICV_9 $T=1062680 598200 1 0 $X=1062680 $Y=592780
X4084 5896 5771 2 1 5902 5897 5868 5755 5878 5848 5872 1233 ICV_9 $T=1063300 628440 0 0 $X=1063300 $Y=628060
X4085 5900 5763 2 1 5922 1127 5720 5744 5864 1136 5884 1233 ICV_9 $T=1063920 567960 0 0 $X=1063920 $Y=567580
X4086 6050 5774 2 1 6092 6005 5680 5994 6044 5993 6021 1233 ICV_9 $T=1096160 588120 0 0 $X=1096160 $Y=587740
X4087 6090 5794 2 1 6114 6101 5935 6016 6030 1163 6080 1233 ICV_9 $T=1099880 557880 1 0 $X=1099880 $Y=552460
X4088 6117 5813 2 1 6141 6140 5829 5682 6027 6098 6106 1233 ICV_9 $T=1103600 699000 0 0 $X=1103600 $Y=698620
X4089 1492 1 2 71 1544 11 1585 49 1233 ICV_11 $T=269080 719160 0 0 $X=269080 $Y=718780
X4090 442 1 2 456 3161 311 3171 3178 1233 ICV_11 $T=563580 699000 0 0 $X=563580 $Y=698620
X4091 526 1 2 3337 3340 311 3354 2931 1233 ICV_11 $T=598920 699000 0 0 $X=598920 $Y=698620
X4092 3327 1 2 3349 3205 553 3353 3430 1233 ICV_11 $T=601400 598200 1 0 $X=601400 $Y=592780
X4093 3451 1 2 3478 3486 3292 3373 3558 1233 ICV_11 $T=624960 648600 1 0 $X=624960 $Y=643180
X4094 599 1 2 3504 3512 3292 3518 3577 1233 ICV_11 $T=628680 658680 0 0 $X=628680 $Y=658300
X4095 3522 1 2 3549 3555 553 3575 3622 1233 ICV_11 $T=635500 588120 0 0 $X=635500 $Y=587740
X4096 3552 1 2 3570 3574 3292 3575 3569 1233 ICV_11 $T=640460 608280 0 0 $X=640460 $Y=607900
X4097 3672 1 2 3711 3712 3292 3750 3194 1233 ICV_11 $T=662780 618360 1 0 $X=662780 $Y=612940
X4098 3790 1 2 3759 3851 3292 3900 3886 1233 ICV_11 $T=691920 658680 1 0 $X=691920 $Y=653260
X4099 3837 1 2 3866 3871 569 3803 3102 1233 ICV_11 $T=692540 699000 1 0 $X=692540 $Y=693580
X4100 3906 1 2 3925 3928 3292 3806 3950 1233 ICV_11 $T=707420 618360 0 0 $X=707420 $Y=617980
X4101 4036 1 2 4065 4097 724 4133 4139 1233 ICV_11 $T=739660 668760 1 0 $X=739660 $Y=663340
X4102 4191 1 2 4209 4200 742 4225 4093 1233 ICV_11 $T=761980 618360 1 0 $X=761980 $Y=612940
X4103 797 1 2 4268 4275 742 811 4270 1233 ICV_11 $T=773760 547800 1 0 $X=773760 $Y=542380
X4104 4296 1 2 4317 4340 724 4217 3370 1233 ICV_11 $T=785540 658680 0 0 $X=785540 $Y=658300
X4105 4291 1 2 4338 4328 742 4304 4353 1233 ICV_11 $T=786160 628440 1 0 $X=786160 $Y=623020
X4106 4506 1 2 4541 4545 839 4595 4619 1233 ICV_11 $T=823980 618360 0 0 $X=823980 $Y=617980
X4107 4509 1 2 4543 4552 837 4481 4572 1233 ICV_11 $T=824600 678840 0 0 $X=824600 $Y=678460
X4108 4787 1 2 4817 4838 839 934 4916 1233 ICV_11 $T=874200 547800 1 0 $X=874200 $Y=542380
X4109 4882 1 2 4926 4938 837 4913 4987 1233 ICV_11 $T=890940 648600 0 0 $X=890940 $Y=648220
X4110 4962 1 2 4984 5000 837 4902 5034 1233 ICV_11 $T=901480 658680 0 0 $X=901480 $Y=658300
X4111 5040 1 2 5050 5067 4818 5082 5060 1233 ICV_11 $T=912640 608280 1 0 $X=912640 $Y=602860
X4112 5187 1 2 5188 5220 4818 5271 1010 1233 ICV_11 $T=938680 608280 0 0 $X=938680 $Y=607900
X4113 5258 1 2 5299 5323 4818 5277 1005 1233 ICV_11 $T=957900 648600 0 0 $X=957900 $Y=648220
X4114 5515 1 2 5505 5595 5560 5584 5585 1233 ICV_11 $T=1008120 618360 0 0 $X=1008120 $Y=617980
X4115 5663 1 2 5691 5695 1025 5702 5663 1233 ICV_11 $T=1024240 588120 1 0 $X=1024240 $Y=582700
X4116 5679 1 2 5697 5707 1025 1117 1106 1233 ICV_11 $T=1026720 547800 1 0 $X=1026720 $Y=542380
X4117 5759 1 2 5786 5805 5560 5765 5811 1233 ICV_11 $T=1045940 638520 1 0 $X=1045940 $Y=633100
X4118 5768 1 2 5791 5815 1121 5822 5824 1233 ICV_11 $T=1047180 557880 1 0 $X=1047180 $Y=552460
X4119 1455 1 2 60 48 53 1233 ICV_14 $T=258540 719160 1 0 $X=258540 $Y=713740
X4120 2410 1 2 259 2359 2459 1233 ICV_14 $T=441440 557880 0 0 $X=441440 $Y=557500
X4121 3406 1 2 3424 3380 3408 1233 ICV_14 $T=611320 608280 0 0 $X=611320 $Y=607900
X4122 737 1 2 747 730 738 1233 ICV_14 $T=730980 547800 1 0 $X=730980 $Y=542380
X4123 3966 1 2 740 731 741 1233 ICV_14 $T=730980 709080 1 0 $X=730980 $Y=703660
X4124 3792 1 2 4075 4045 4073 1233 ICV_14 $T=735940 567960 0 0 $X=735940 $Y=567580
X4125 3914 1 2 4070 4093 4123 1233 ICV_14 $T=745240 608280 1 0 $X=745240 $Y=602860
X4126 4691 1 2 4710 877 4723 1233 ICV_14 $T=859940 719160 1 0 $X=859940 $Y=713740
X4127 4688 1 2 4633 4425 4488 1233 ICV_14 $T=868620 628440 0 0 $X=868620 $Y=628060
X4128 4701 1 2 4880 4834 4868 1233 ICV_14 $T=878540 688920 1 0 $X=878540 $Y=683500
X4129 4790 1 2 4897 4845 4833 1233 ICV_14 $T=880400 648600 1 0 $X=880400 $Y=643180
X4130 4725 1 2 4930 935 937 1233 ICV_14 $T=887220 699000 0 0 $X=887220 $Y=698620
X4131 4893 1 2 4886 4885 4906 1233 ICV_14 $T=888460 678840 1 0 $X=888460 $Y=673420
X4132 891 1 2 4943 4914 4904 1233 ICV_14 $T=890940 598200 1 0 $X=890940 $Y=592780
X4133 4759 1 2 5080 5113 5143 1233 ICV_14 $T=926280 688920 1 0 $X=926280 $Y=683500
X4134 5184 1 2 5191 5116 5147 1233 ICV_14 $T=932480 678840 0 0 $X=932480 $Y=678460
X4135 5199 1 2 5264 5203 5216 1233 ICV_14 $T=943640 608280 1 0 $X=943640 $Y=602860
X4136 5407 1 2 5443 5410 5436 1233 ICV_14 $T=983320 567960 1 0 $X=983320 $Y=562540
X4137 1045 1 2 1076 5454 5488 1233 ICV_14 $T=990140 628440 1 0 $X=990140 $Y=623020
X4138 5634 1 2 5649 5594 5571 1233 ICV_14 $T=1013700 668760 1 0 $X=1013700 $Y=663340
X4139 5671 1 2 1117 5665 5728 1233 ICV_14 $T=1032920 547800 0 0 $X=1032920 $Y=547420
X4140 5518 1 2 5512 5667 5714 1233 ICV_14 $T=1032920 638520 1 0 $X=1032920 $Y=633100
X4141 5638 1 2 5778 5743 5769 1233 ICV_14 $T=1039740 557880 0 0 $X=1039740 $Y=557500
X4142 5590 1 2 5812 5737 5784 1233 ICV_14 $T=1045320 678840 1 0 $X=1045320 $Y=673420
X4143 6133 1 2 6089 6105 6099 1233 ICV_14 $T=1105460 658680 1 0 $X=1105460 $Y=653260
X4144 1484 2 1524 1 1524 70 1233 ICV_16 $T=272180 699000 0 0 $X=272180 $Y=698620
X4145 1765 2 1785 1 1681 1543 1233 ICV_16 $T=318060 688920 0 0 $X=318060 $Y=688540
X4146 2425 2 2414 1 2219 2432 1233 ICV_16 $T=437100 648600 0 0 $X=437100 $Y=648220
X4147 2401 2 2501 1 2501 2474 1233 ICV_16 $T=449500 648600 1 0 $X=449500 $Y=643180
X4148 3004 2 3166 1 3166 3125 1233 ICV_16 $T=568540 638520 1 0 $X=568540 $Y=633100
X4149 626 2 3562 1 3513 3503 1233 ICV_16 $T=641700 709080 1 0 $X=641700 $Y=703660
X4150 3707 2 3755 1 3707 672 1233 ICV_16 $T=675800 557880 1 0 $X=675800 $Y=552460
X4151 4145 2 787 1 4013 4208 1233 ICV_16 $T=763220 699000 0 0 $X=763220 $Y=698620
X4152 4357 2 4293 1 4293 818 1233 ICV_16 $T=795460 578040 0 0 $X=795460 $Y=577660
X4153 4082 2 836 1 4082 4464 1233 ICV_16 $T=814060 719160 1 0 $X=814060 $Y=713740
X4154 4752 2 4757 1 4477 4752 1233 ICV_16 $T=863660 648600 1 0 $X=863660 $Y=643180
X4155 4594 2 4905 1 4929 4942 1233 ICV_16 $T=894660 588120 0 0 $X=894660 $Y=587740
X4156 990 2 5139 1 5139 5170 1233 ICV_16 $T=934340 588120 0 0 $X=934340 $Y=587740
X4157 5504 2 5539 1 4878 5456 1233 ICV_16 $T=1003160 588120 0 0 $X=1003160 $Y=587740
X4158 5566 2 5568 1 5566 1087 1233 ICV_16 $T=1008120 578040 1 0 $X=1008120 $Y=572620
X4159 5417 2 5582 1 5417 5590 1233 ICV_16 $T=1010600 678840 0 0 $X=1010600 $Y=678460
X4160 5575 2 5659 1 5659 5671 1233 ICV_16 $T=1023620 578040 1 0 $X=1023620 $Y=572620
X4161 5925 2 5932 1 5925 5937 1233 ICV_16 $T=1073220 578040 0 0 $X=1073220 $Y=577660
X4162 5937 2 6146 1 6146 1172 1233 ICV_16 $T=1111040 547800 1 0 $X=1111040 $Y=542380
X4163 220 1960 1 2 INV6CK $T=409820 608280 0 180 $X=404240 $Y=602860
X4164 2270 220 1 2 INV6CK $T=412300 578040 0 0 $X=412300 $Y=577660
X4165 3860 2270 1 2 INV6CK $T=696260 578040 0 0 $X=696260 $Y=577660
X4166 4327 815 1 2 INV6CK $T=788640 578040 0 0 $X=788640 $Y=577660
X4167 982 5425 1 2 INV6CK $T=987040 547800 0 180 $X=981460 $Y=542380
X4168 5849 5825 5827 5840 4441 1 2 AN4 $T=1059580 678840 0 180 $X=1053380 $Y=673420
X4169 1323 1348 1336 1 2 ND2 $T=238700 567960 0 180 $X=236840 $Y=562540
X4170 1278 1354 1317 1 2 ND2 $T=242420 547800 1 0 $X=242420 $Y=542380
X4171 89 96 1633 1 2 ND2 $T=293880 567960 0 180 $X=292020 $Y=562540
X4172 1741 1745 1766 1 2 ND2 $T=313100 598200 1 0 $X=313100 $Y=592780
X4173 1762 1737 1772 1 2 ND2 $T=314960 598200 0 0 $X=314960 $Y=597820
X4174 2256 2380 2386 1 2 ND2 $T=428420 578040 1 0 $X=428420 $Y=572620
X4175 2687 2583 2728 1 2 ND2 $T=489180 598200 1 0 $X=489180 $Y=592780
X4176 2775 2790 2825 1 2 ND2 $T=505300 598200 0 0 $X=505300 $Y=597820
X4177 3177 3181 3189 1 2 ND2 $T=572260 668760 1 0 $X=572260 $Y=663340
X4178 3177 3195 2970 1 2 ND2 $T=574120 668760 1 0 $X=574120 $Y=663340
X4179 3189 3211 2970 1 2 ND2 $T=580940 668760 1 0 $X=580940 $Y=663340
X4180 3241 3288 3269 1 2 ND2 $T=593960 658680 1 0 $X=593960 $Y=653260
X4181 3339 3360 3303 1 2 ND2 $T=608220 628440 1 180 $X=606360 $Y=628060
X4182 3527 3243 3494 1 2 ND2 $T=638600 699000 1 0 $X=638600 $Y=693580
X4183 3533 3579 3494 1 2 ND2 $T=649140 699000 0 180 $X=647280 $Y=693580
X4184 3608 645 3633 1 2 ND2 $T=654100 537720 0 0 $X=654100 $Y=537340
X4185 606 3633 641 1 2 ND2 $T=655960 537720 0 0 $X=655960 $Y=537340
X4186 5535 5542 5466 1 2 ND2 $T=1003780 658680 1 0 $X=1003780 $Y=653260
X4187 4281 804 1 2 INV8CK $T=779340 709080 0 0 $X=779340 $Y=708700
X4188 3860 4327 1 2 INV8CK $T=788640 588120 0 0 $X=788640 $Y=587740
X4189 4327 4281 1 2 INV8CK $T=788640 709080 0 0 $X=788640 $Y=708700
X4190 5425 5370 1 2 INV8CK $T=991380 547800 0 0 $X=991380 $Y=547420
X4191 3303 3306 2 3339 3351 3306 1 AOI22HP $T=597060 638520 1 0 $X=597060 $Y=633100
X4192 3406 3444 2 3384 3502 3444 1 AOI22HP $T=623100 628440 1 0 $X=623100 $Y=623020
X4193 1317 1318 2 1278 1346 1318 1 AOI22H $T=233740 547800 1 0 $X=233740 $Y=542380
X4194 1336 1352 2 1323 1351 1352 1 AOI22H $T=247380 567960 0 180 $X=239940 $Y=562540
X4195 3195 3216 3181 3211 1 2 ND3P $T=575980 668760 1 0 $X=575980 $Y=663340
X4196 843 2 786 1 4477 NR2P $T=819020 638520 1 180 $X=815300 $Y=638140
X4197 778 2 843 1 4500 NR2P $T=819640 648600 1 0 $X=819640 $Y=643180
X4198 1048 2 1038 1 5403 NR2P $T=985180 688920 0 0 $X=985180 $Y=688540
X4199 880 2 1053 1 5422 NR2P $T=987040 678840 1 0 $X=987040 $Y=673420
X4200 1308 2 1334 1326 1316 1 1274 FA1S $T=236840 648600 0 180 $X=225060 $Y=643180
X4201 1299 2 1364 1347 1353 1 1311 FA1S $T=244280 668760 0 180 $X=232500 $Y=663340
X4202 1293 2 1355 1379 1320 1 1309 FA1S $T=244900 678840 1 180 $X=233120 $Y=678460
X4203 1353 2 1378 1368 1360 1 1320 FA1S $T=246140 688920 1 180 $X=234360 $Y=688540
X4204 1349 2 1366 1330 1358 1 1292 FA1S $T=246760 628440 1 180 $X=234980 $Y=628060
X4205 1357 2 1382 1371 1363 1 1330 FA1S $T=247380 618360 1 180 $X=235600 $Y=617980
X4206 1358 2 1394 1341 1367 1 1326 FA1S $T=247380 638520 1 180 $X=235600 $Y=638140
X4207 1336 2 1401 1374 1356 1 1289 FA1S $T=248000 578040 1 180 $X=236220 $Y=577660
X4208 1359 2 20 1392 1365 1 1335 FA1S $T=248000 648600 1 180 $X=236220 $Y=648220
X4209 1356 2 3 1377 1389 1 1395 FA1S $T=237460 588120 1 0 $X=237460 $Y=582700
X4210 1334 2 1391 1383 1359 1 1342 FA1S $T=249240 648600 0 180 $X=237460 $Y=643180
X4211 36 2 14 1386 1361 1 1318 FA1S $T=249860 547800 1 180 $X=238080 $Y=547420
X4212 1325 2 1402 1405 1381 1 1273 FA1S $T=249860 598200 1 180 $X=238080 $Y=597820
X4213 1269 2 1370 1406 1357 1 1344 FA1S $T=249860 608280 1 180 $X=238080 $Y=607900
X4214 1316 2 1411 1419 1342 1 1347 FA1S $T=250480 658680 1 180 $X=238700 $Y=658300
X4215 1371 2 22 1416 1385 1 1341 FA1S $T=251100 638520 0 180 $X=239320 $Y=633100
X4216 1364 2 1426 1412 1335 1 1355 FA1S $T=252960 668760 1 180 $X=241180 $Y=668380
X4217 1379 2 1362 1420 1390 1 1435 FA1S $T=242420 678840 1 0 $X=242420 $Y=673420
X4218 1402 2 4 1431 1436 1 1370 FA1S $T=256680 608280 0 180 $X=244900 $Y=602860
X4219 1411 2 1448 1442 1433 1 1368 FA1S $T=256680 668760 0 180 $X=244900 $Y=663340
X4220 1378 2 1457 1459 1429 1 1362 FA1S $T=256680 688920 0 180 $X=244900 $Y=683500
X4221 1423 2 5 49 1439 1 1374 FA1S $T=257920 578040 0 180 $X=246140 $Y=572620
X4222 1317 2 6 1450 1423 1 1352 FA1S $T=258540 567960 1 180 $X=246760 $Y=567580
X4223 1360 2 1400 1477 1453 1 1390 FA1S $T=259780 688920 1 180 $X=248000 $Y=688540
X4224 1452 2 1473 1458 1440 1 1363 FA1S $T=261020 628440 0 180 $X=249240 $Y=623020
X4225 1381 2 1466 1463 1452 1 1406 FA1S $T=262260 618360 0 180 $X=250480 $Y=612940
X4226 1463 2 9 56 1468 1 1382 FA1S $T=262880 618360 1 180 $X=251100 $Y=617980
X4227 1366 2 1446 1432 1494 1 1367 FA1S $T=253580 638520 0 0 $X=253580 $Y=638140
X4228 1394 2 1447 1451 1472 1 1419 FA1S $T=253580 658680 0 0 $X=253580 $Y=658300
X4229 1313 2 1489 1395 1482 1 1322 FA1S $T=265980 588120 1 180 $X=254200 $Y=587740
X4230 1482 2 1498 1493 1488 1 1405 FA1S $T=267840 598200 0 180 $X=256060 $Y=592780
X4231 1489 2 8 65 1471 1 1488 FA1S $T=259780 598200 0 0 $X=259780 $Y=597820
X4232 1494 2 15 1547 1470 1 1383 FA1S $T=271560 648600 0 180 $X=259780 $Y=643180
X4233 1412 2 1475 1474 1478 1 1532 FA1S $T=261020 668760 0 0 $X=261020 $Y=668380
X4234 1294 2 1532 1499 1435 1 1522 FA1S $T=263500 678840 1 0 $X=263500 $Y=673420
X4235 1453 2 1495 1516 1538 1 1567 FA1S $T=267220 699000 1 0 $X=267220 $Y=693580
X4236 1420 2 1555 1581 1523 1 1570 FA1S $T=271560 688920 1 0 $X=271560 $Y=683500
X4237 1521 2 1650 1621 1541 1 1549 FA1S $T=287060 658680 0 180 $X=275280 $Y=653260
X4238 1597 2 1615 1610 1603 1 1541 FA1S $T=288300 668760 1 180 $X=276520 $Y=668380
X4239 1527 2 1626 1597 1609 1 1526 FA1S $T=288920 668760 0 180 $X=277140 $Y=663340
X4240 1499 2 1605 1570 1567 1 1609 FA1S $T=277760 678840 1 0 $X=277760 $Y=673420
X4241 1605 2 1573 1594 1586 1 1603 FA1S $T=280860 688920 0 0 $X=280860 $Y=688540
X4242 1621 2 1639 1647 1624 1 1575 FA1S $T=293260 658680 1 180 $X=281480 $Y=658300
X4243 1614 2 1643 1632 1673 1 1622 FA1S $T=300700 608280 1 180 $X=288920 $Y=607900
X4244 1608 2 1676 1728 1575 1 1618 FA1S $T=301320 648600 0 180 $X=289540 $Y=643180
X4245 1670 2 1691 1694 1663 1 1632 FA1S $T=302560 618360 1 180 $X=290780 $Y=617980
X4246 1619 2 1637 1670 1680 1 1607 FA1S $T=302560 628440 1 180 $X=290780 $Y=628060
X4247 1626 2 1630 1640 1660 1 1610 FA1S $T=290780 678840 1 0 $X=290780 $Y=673420
X4248 1676 2 1693 1686 1666 1 1637 FA1S $T=303800 638520 0 180 $X=292020 $Y=633100
X4249 1624 2 1678 1667 1699 1 1680 FA1S $T=297600 658680 0 0 $X=297600 $Y=658300
X4250 107 2 1665 1719 1677 1 115 FA1S $T=298220 537720 0 0 $X=298220 $Y=537340
X4251 1650 2 1671 1709 1674 1 1728 FA1S $T=298220 648600 0 0 $X=298220 $Y=648220
X4252 1673 2 1754 1746 1736 1 1679 FA1S $T=314340 608280 1 180 $X=302560 $Y=607900
X4253 1735 2 1718 1634 1748 1 129 FA1S $T=306280 688920 0 0 $X=306280 $Y=688540
X4254 119 2 1716 1547 1749 1 130 FA1S $T=306280 699000 0 0 $X=306280 $Y=698620
X4255 1749 2 1711 1485 1735 1 133 FA1S $T=308140 699000 1 0 $X=308140 $Y=693580
X4256 1768 2 1547 125 1774 1 1793 FA1S $T=311240 648600 1 0 $X=311240 $Y=643180
X4257 1774 2 1485 124 1813 1 1812 FA1S $T=311860 658680 0 0 $X=311860 $Y=658300
X4258 134 2 1747 1504 1800 1 140 FA1S $T=316200 537720 0 0 $X=316200 $Y=537340
X4259 1820 2 56 141 1768 1 1843 FA1S $T=321160 638520 0 0 $X=321160 $Y=638140
X4260 1838 2 145 1814 143 1 135 FA1S $T=334800 719160 1 180 $X=323020 $Y=718780
X4261 1845 2 1857 1865 1850 1 1814 FA1S $T=336040 709080 0 180 $X=324260 $Y=703660
X4262 1813 2 1634 138 1868 1 1860 FA1S $T=325500 658680 0 0 $X=325500 $Y=658300
X4263 1762 2 1833 1832 1830 1 1784 FA1S $T=337900 608280 0 180 $X=326120 $Y=602860
X4264 150 2 1862 1893 151 1 142 FA1S $T=342240 537720 1 180 $X=330460 $Y=537340
X4265 1868 2 1740 152 1874 1 1903 FA1S $T=332940 648600 1 0 $X=332940 $Y=643180
X4266 1874 2 1681 157 1867 1 1914 FA1S $T=334180 638520 0 0 $X=334180 $Y=638140
X4267 6186 2 1845 1900 1838 1 144 FA1S $T=345960 709080 1 180 $X=334180 $Y=708700
X4268 6187 2 1965 1897 1884 1 1859 FA1S $T=347200 699000 1 180 $X=335420 $Y=698620
X4269 1897 2 1938 1910 1890 1 1865 FA1S $T=348440 709080 0 180 $X=336660 $Y=703660
X4270 1857 2 1910 158 1907 1 147 FA1S $T=348440 719160 1 180 $X=336660 $Y=718780
X4271 1889 2 65 159 1820 1 1926 FA1S $T=337280 638520 1 0 $X=337280 $Y=633100
X4272 156 2 1901 1846 1949 1 164 FA1S $T=339140 557880 0 0 $X=339140 $Y=557500
X4273 1867 2 1844 165 1964 1 1895 FA1S $T=357740 618360 1 180 $X=345960 $Y=617980
X4274 6188 2 1947 1910 1938 1 1884 FA1S $T=347200 709080 0 0 $X=347200 $Y=708700
X4275 6189 2 1976 2001 1859 1 1900 FA1S $T=362080 699000 0 180 $X=350300 $Y=693580
X4276 1976 2 2034 1990 1980 1 1850 FA1S $T=362700 709080 0 180 $X=350920 $Y=703660
X4277 1949 2 1962 1856 1958 1 184 FA1S $T=353400 557880 0 0 $X=353400 $Y=557500
X4278 1990 2 2011 173 2003 1 169 FA1S $T=366420 719160 0 180 $X=354640 $Y=713740
X4279 6190 2 2021 2029 2000 1 1965 FA1S $T=367040 688920 1 180 $X=355260 $Y=688540
X4280 1890 2 185 189 2005 1 1907 FA1S $T=367040 719160 1 180 $X=355260 $Y=718780
X4281 6191 2 2064 2068 2046 1 2001 FA1S $T=375100 699000 0 180 $X=363320 $Y=693580
X4282 2046 2 2024 2060 2038 1 1980 FA1S $T=376340 699000 1 180 $X=364560 $Y=698620
X4283 2060 2 193 2075 2069 1 2003 FA1S $T=378200 719160 0 180 $X=366420 $Y=713740
X4284 2064 2 2086 2076 2084 1 2034 FA1S $T=381920 709080 1 180 $X=370140 $Y=708700
X4285 2076 2 195 2102 2085 1 2005 FA1S $T=381920 719160 1 180 $X=370140 $Y=718780
X4286 2029 2 2105 2099 2092 1 2038 FA1S $T=383160 688920 1 180 $X=371380 $Y=688540
X4287 2090 2 1386 196 2094 1 2128 FA1S $T=375100 578040 0 0 $X=375100 $Y=577660
X4288 2094 2 49 201 1889 1 2132 FA1S $T=375720 598200 1 0 $X=375720 $Y=592780
X4289 194 2 2047 1912 2103 1 206 FA1S $T=376340 547800 1 0 $X=376340 $Y=542380
X4290 6192 2 2080 2155 2113 1 2068 FA1S $T=389980 699000 1 180 $X=378200 $Y=698620
X4291 6193 2 2178 2159 2141 1 2000 FA1S $T=396180 688920 1 180 $X=384400 $Y=688540
X4292 2155 2 2160 2125 2165 1 2084 FA1S $T=396180 709080 0 180 $X=384400 $Y=703660
X4293 6194 2 2175 2168 2174 1 2113 FA1S $T=396800 699000 0 180 $X=385020 $Y=693580
X4294 2161 2 2189 2137 2048 1 2206 FA1S $T=388120 547800 0 0 $X=388120 $Y=547420
X4295 209 2 2176 2022 2122 1 2228 FA1S $T=390600 547800 1 0 $X=390600 $Y=542380
X4296 6195 2 2180 2205 2211 1 2159 FA1S $T=403620 678840 0 180 $X=391840 $Y=673420
X4297 2085 2 2201 2152 2213 1 217 FA1S $T=395560 719160 0 0 $X=395560 $Y=718780
X4298 2174 2 2187 2199 2203 1 2099 FA1S $T=398040 688920 0 0 $X=398040 $Y=688540
X4299 2165 2 2200 2214 2197 1 2075 FA1S $T=399280 709080 1 0 $X=399280 $Y=703660
X4300 2286 2 2263 2262 2319 1 2352 FA1S $T=411060 567960 1 0 $X=411060 $Y=562540
X4301 2318 2 2337 2297 2324 1 241 FA1S $T=415400 699000 0 0 $X=415400 $Y=698620
X4302 2368 2 2361 2336 2302 1 2411 FA1S $T=422840 547800 0 0 $X=422840 $Y=547420
X4303 240 2 2340 2323 2348 1 244 FA1S $T=422840 719160 0 0 $X=422840 $Y=718780
X4304 2381 2 2343 2311 2367 1 2422 FA1S $T=424700 688920 1 0 $X=424700 $Y=683500
X4305 2394 2 2344 2339 2326 1 248 FA1S $T=426560 709080 1 0 $X=426560 $Y=703660
X4306 243 2 2332 239 2261 1 2433 FA1S $T=427180 547800 1 0 $X=427180 $Y=542380
X4307 2392 2 2364 2371 2381 1 2429 FA1S $T=427180 688920 0 0 $X=427180 $Y=688540
X4308 2398 2 2281 2382 2318 1 2458 FA1S $T=427800 699000 0 0 $X=427800 $Y=698620
X4309 2403 2 2378 2354 2455 1 2456 FA1S $T=429660 668760 1 0 $X=429660 $Y=663340
X4310 6196 2 2379 2392 2448 1 2457 FA1S $T=429660 678840 0 0 $X=429660 $Y=678460
X4311 6197 2 2384 2377 2403 1 2448 FA1S $T=430280 678840 1 0 $X=430280 $Y=673420
X4312 2464 2 2374 2417 2394 1 2503 FA1S $T=438960 709080 0 0 $X=438960 $Y=708700
X4313 2467 2 2434 2398 2429 1 2509 FA1S $T=439580 699000 1 0 $X=439580 $Y=693580
X4314 2468 2 2443 252 2503 1 262 FA1S $T=439580 719160 0 0 $X=439580 $Y=718780
X4315 2475 2 2437 2464 2458 1 267 FA1S $T=440820 709080 1 0 $X=440820 $Y=703660
X4316 2498 2 2480 2456 2452 1 2527 FA1S $T=445160 668760 0 0 $X=445160 $Y=668380
X4317 2499 2 2471 2422 2488 1 2536 FA1S $T=445160 688920 0 0 $X=445160 $Y=688540
X4318 2502 2 2527 2477 2475 1 2542 FA1S $T=445780 678840 0 0 $X=445780 $Y=678460
X4319 6198 2 2476 2532 2463 1 2569 FA1S $T=446400 658680 0 0 $X=446400 $Y=658300
X4320 6199 2 2563 2553 2548 1 261 FA1S $T=460660 537720 1 180 $X=448880 $Y=537340
X4321 6200 2 2537 2595 2582 1 2524 FA1S $T=466860 557880 0 180 $X=455080 $Y=552460
X4322 2559 2 2509 2534 269 1 2602 FA1S $T=455080 719160 1 0 $X=455080 $Y=713740
X4323 6201 2 2549 2498 2554 1 2600 FA1S $T=457560 668760 1 0 $X=457560 $Y=663340
X4324 6202 2 2550 2600 2502 1 2637 FA1S $T=457560 678840 1 0 $X=457560 $Y=673420
X4325 6203 2 2522 2601 2559 1 2615 FA1S $T=457560 709080 1 0 $X=457560 $Y=703660
X4326 2581 2 2551 2499 2552 1 2628 FA1S $T=458800 688920 0 0 $X=458800 $Y=688540
X4327 6204 2 2569 2533 2467 1 2601 FA1S $T=458800 699000 1 0 $X=458800 $Y=693580
X4328 6205 2 2616 2567 2580 1 2640 FA1S $T=460040 588120 1 0 $X=460040 $Y=582700
X4329 6206 2 2568 2579 2590 1 2532 FA1S $T=461900 658680 0 0 $X=461900 $Y=658300
X4330 2618 2 2652 2650 2626 1 272 FA1S $T=474920 668760 1 180 $X=463140 $Y=668380
X4331 2604 2 2536 2529 2468 1 289 FA1S $T=463140 709080 0 0 $X=463140 $Y=708700
X4332 6207 2 2457 2511 2581 1 2653 FA1S $T=465000 688920 1 0 $X=465000 $Y=683500
X4333 6208 2 2608 2594 2631 1 2692 FA1S $T=466240 567960 0 0 $X=466240 $Y=567580
X4334 2627 2 2542 290 2602 1 296 FA1S $T=466860 719160 1 0 $X=466860 $Y=713740
X4335 2656 2 2684 2670 2625 1 6209 FA1S $T=481740 638520 0 180 $X=469960 $Y=633100
X4336 2657 2 2673 2691 2618 1 278 FA1S $T=481740 678840 1 180 $X=469960 $Y=678460
X4337 6210 2 2679 2694 2666 1 2621 FA1S $T=482360 578040 1 180 $X=470580 $Y=577660
X4338 2626 2 2677 2635 2656 1 6211 FA1S $T=482360 668760 0 180 $X=470580 $Y=663340
X4339 6212 2 2653 2645 2637 1 2690 FA1S $T=472440 688920 0 0 $X=472440 $Y=688540
X4340 2645 2 2629 2628 2604 1 308 FA1S $T=473060 699000 1 0 $X=473060 $Y=693580
X4341 6213 2 2627 2615 2690 1 309 FA1S $T=473060 709080 1 0 $X=473060 $Y=703660
X4342 2693 2 2720 2724 2685 1 2650 FA1S $T=489180 678840 0 180 $X=477400 $Y=673420
X4343 6214 2 302 2674 2682 1 319 FA1S $T=479880 547800 1 0 $X=479880 $Y=542380
X4344 6215 2 2695 2675 2706 1 2768 FA1S $T=483600 547800 0 0 $X=483600 $Y=547420
X4345 2730 2 2763 2751 2693 1 2691 FA1S $T=495380 678840 1 180 $X=483600 $Y=678460
X4346 2731 2 2771 2777 2714 1 2689 FA1S $T=495380 688920 0 180 $X=483600 $Y=683500
X4347 6216 2 2755 2769 2700 1 2694 FA1S $T=496000 578040 1 180 $X=484220 $Y=577660
X4348 2716 2 2730 2689 2657 1 325 FA1S $T=485460 699000 1 0 $X=485460 $Y=693580
X4349 2759 2 2731 2778 2716 1 313 FA1S $T=499100 699000 1 180 $X=487320 $Y=698620
X4350 6217 2 2772 2733 2765 1 2797 FA1S $T=492280 588120 1 0 $X=492280 $Y=582700
X4351 6218 2 2732 2792 2748 1 2816 FA1S $T=493520 557880 1 0 $X=493520 $Y=552460
X4352 2813 2 2828 2740 2822 1 2778 FA1S $T=509640 688920 0 180 $X=497860 $Y=683500
X4353 2823 2 2813 2838 2759 1 329 FA1S $T=510880 699000 0 180 $X=499100 $Y=693580
X4354 2832 2 2808 2855 2704 1 2866 FA1S $T=503440 618360 1 0 $X=503440 $Y=612940
X4355 6219 2 2872 2854 2837 1 2800 FA1S $T=515840 588120 0 180 $X=504060 $Y=582700
X4356 2859 2 2978 2852 2866 1 2826 FA1S $T=518320 618360 1 180 $X=506540 $Y=617980
X4357 2860 2 2859 2892 2867 1 341 FA1S $T=518320 638520 0 180 $X=506540 $Y=633100
X4358 6220 2 2850 2815 2836 1 2865 FA1S $T=507160 567960 0 0 $X=507160 $Y=567580
X4359 2844 2 2881 2842 2804 1 2897 FA1S $T=507780 608280 0 0 $X=507780 $Y=607900
X4360 2852 2 2809 2882 2747 1 2911 FA1S $T=507780 628440 0 0 $X=507780 $Y=628060
X4361 2867 2 2891 2826 2861 1 347 FA1S $T=519560 638520 1 180 $X=507780 $Y=638140
X4362 6221 2 2847 2841 2879 1 2863 FA1S $T=510260 588120 0 0 $X=510260 $Y=587740
X4363 6222 2 2898 2844 2736 1 2922 FA1S $T=510260 598200 0 0 $X=510260 $Y=597820
X4364 2873 2 2760 2900 2906 1 2916 FA1S $T=510880 648600 0 0 $X=510880 $Y=648220
X4365 2861 2 2873 2907 2899 1 352 FA1S $T=523280 658680 0 180 $X=511500 $Y=653260
X4366 2878 2 2909 2754 2853 1 2913 FA1S $T=511500 688920 1 0 $X=511500 $Y=683500
X4367 2888 2 2928 2913 2823 1 355 FA1S $T=523280 699000 0 180 $X=511500 $Y=693580
X4368 2862 2 2930 2840 2908 1 2853 FA1S $T=523900 668760 0 180 $X=512120 $Y=663340
X4369 2896 2 2878 2919 2888 1 358 FA1S $T=523900 688920 1 180 $X=512120 $Y=688540
X4370 2884 2 2753 2862 2871 1 2919 FA1S $T=512740 668760 0 0 $X=512740 $Y=668380
X4371 2899 2 2884 2916 2896 1 353 FA1S $T=524520 678840 0 180 $X=512740 $Y=673420
X4372 6223 2 2816 2880 2939 1 2941 FA1S $T=515840 557880 1 0 $X=515840 $Y=552460
X4373 6224 2 2929 2890 2893 1 2939 FA1S $T=517700 547800 0 0 $X=517700 $Y=547420
X4374 6225 2 2827 2903 2926 1 2960 FA1S $T=518320 567960 1 0 $X=518320 $Y=562540
X4375 2891 2 2902 2946 2911 1 2907 FA1S $T=520180 638520 1 0 $X=520180 $Y=633100
X4376 2855 2 2968 2974 2957 1 2902 FA1S $T=532580 628440 1 180 $X=520800 $Y=628060
X4377 2946 2 2963 2820 2954 1 2906 FA1S $T=532580 648600 0 180 $X=520800 $Y=643180
X4378 2904 2 2897 2832 2944 1 2892 FA1S $T=521420 608280 0 0 $X=521420 $Y=607900
X4379 2900 2 2975 2833 2918 1 2871 FA1S $T=533200 658680 1 180 $X=521420 $Y=658300
X4380 6226 2 2921 2935 2910 1 2966 FA1S $T=523280 588120 1 0 $X=523280 $Y=582700
X4381 6227 2 2927 2973 2803 1 2990 FA1S $T=523900 598200 1 0 $X=523900 $Y=592780
X4382 6228 2 2990 2982 2922 1 2895 FA1S $T=536300 598200 1 180 $X=524520 $Y=597820
X4383 2963 2 2992 3000 2979 1 2918 FA1S $T=536300 648600 1 180 $X=524520 $Y=648220
X4384 2909 2 3008 2987 2848 1 2933 FA1S $T=536920 668760 0 180 $X=525140 $Y=663340
X4385 2928 2 2980 2739 2933 1 2838 FA1S $T=525760 688920 1 0 $X=525760 $Y=683500
X4386 2980 2 3022 3002 2993 1 2822 FA1S $T=538780 678840 1 180 $X=527000 $Y=678460
X4387 2982 2 3015 3030 2717 1 2944 FA1S $T=539400 608280 0 180 $X=527620 $Y=602860
X4388 6229 2 2938 2961 2952 1 3009 FA1S $T=528860 578040 1 0 $X=528860 $Y=572620
X4389 3030 2 3047 2998 3050 1 2978 FA1S $T=549320 608280 1 180 $X=537540 $Y=607900
X4390 3043 2 3044 3127 3054 1 3007 FA1S $T=549940 588120 1 180 $X=538160 $Y=587740
X4391 2973 2 3043 3062 3055 1 3015 FA1S $T=550560 598200 1 180 $X=538780 $Y=597820
X4392 3047 2 3078 3066 3056 1 2957 FA1S $T=551180 618360 0 180 $X=539400 $Y=612940
X4393 2993 2 3072 3045 3027 1 2777 FA1S $T=551180 688920 0 180 $X=539400 $Y=683500
X4394 2882 2 3090 2995 3074 1 2954 FA1S $T=553660 638520 1 180 $X=541880 $Y=638140
X4395 6230 2 3088 3039 3071 1 2898 FA1S $T=554280 608280 0 180 $X=542500 $Y=602860
X4396 2842 2 3100 3079 3007 1 3050 FA1S $T=551800 608280 0 0 $X=551800 $Y=607900
X4397 3114 2 3129 3133 3049 1 3084 FA1S $T=564200 578040 1 180 $X=552420 $Y=577660
X4398 3054 2 3111 3143 3118 1 3066 FA1S $T=564200 598200 0 180 $X=552420 $Y=592780
X4399 3088 2 3144 3084 3119 1 3055 FA1S $T=564820 598200 1 180 $X=553040 $Y=597820
X4400 2975 2 3160 3138 3145 1 2908 FA1S $T=567920 658680 1 180 $X=556140 $Y=658300
X4401 6231 2 3169 3115 3137 1 3071 FA1S $T=569780 608280 0 180 $X=558000 $Y=602860
X4402 3145 2 3174 3158 3164 1 2987 FA1S $T=572260 668760 0 180 $X=560480 $Y=663340
X4403 6232 2 3173 3142 3114 1 3137 FA1S $T=567920 578040 0 0 $X=567920 $Y=577660
X4404 3197 2 3198 3179 3162 1 488 FA1S $T=571640 557880 1 0 $X=571640 $Y=552460
X4405 2968 2 3200 3201 3227 1 3074 FA1S $T=585900 638520 0 180 $X=574120 $Y=633100
X4406 3213 2 3223 378 3193 1 3253 FA1S $T=575360 567960 1 0 $X=575360 $Y=562540
X4407 3224 2 3271 3202 3235 1 475 FA1S $T=587760 547800 1 180 $X=575980 $Y=547420
X4408 3227 2 3258 3215 3256 1 3000 FA1S $T=589620 638520 1 180 $X=577840 $Y=638140
X4409 3270 2 3244 3232 3252 1 3274 FA1S $T=584040 557880 0 0 $X=584040 $Y=557500
X4410 3279 2 3247 3267 3280 1 3308 FA1S $T=587140 567960 0 0 $X=587140 $Y=567580
X4411 3287 2 3197 3274 3224 1 530 FA1S $T=589000 547800 0 0 $X=589000 $Y=547420
X4412 3305 2 3313 3276 3300 1 3338 FA1S $T=593340 588120 0 0 $X=593340 $Y=587740
X4413 3385 2 3382 3332 3362 1 3445 FA1S $T=608840 588120 0 0 $X=608840 $Y=587740
X4414 574 2 3376 3381 3375 1 3437 FA1S $T=610700 547800 1 0 $X=610700 $Y=542380
X4415 3398 2 502 3324 3377 1 3425 FA1S $T=610700 567960 0 0 $X=610700 $Y=567580
X4416 3439 2 3352 3411 3446 1 3475 FA1S $T=618140 547800 0 0 $X=618140 $Y=547420
X4417 601 2 3383 3347 3448 1 3520 FA1S $T=624340 567960 0 0 $X=624340 $Y=567580
X4418 3474 2 3437 3419 3439 1 3535 FA1S $T=624960 547800 1 0 $X=624960 $Y=542380
X4419 3525 2 3392 3398 3520 1 3563 FA1S $T=631780 557880 0 0 $X=631780 $Y=557500
X4420 3538 2 3475 3304 3519 1 3580 FA1S $T=634260 557880 1 0 $X=634260 $Y=552460
X4421 1491 1469 1479 2 1 XNR2HS $T=265980 547800 1 180 $X=260400 $Y=547420
X4422 72 74 77 2 1 XNR2HS $T=273420 537720 0 0 $X=273420 $Y=537340
X4423 1551 76 78 2 1 XNR2HS $T=275280 547800 1 0 $X=275280 $Y=542380
X4424 1551 59 82 2 1 XNR2HS $T=283340 537720 0 0 $X=283340 $Y=537340
X4425 1551 1611 86 2 1 XNR2HS $T=285200 547800 1 0 $X=285200 $Y=542380
X4426 1578 1604 87 2 1 XNR2HS $T=285820 557880 1 0 $X=285820 $Y=552460
X4427 1551 1638 1644 2 1 XNR2HS $T=292020 557880 1 0 $X=292020 $Y=552460
X4428 1675 1592 1658 2 1 XNR2HS $T=300080 567960 1 180 $X=294500 $Y=567580
X4429 1675 1616 1672 2 1 XNR2HS $T=302560 567960 0 180 $X=296980 $Y=562540
X4430 1675 1611 1704 2 1 XNR2HS $T=301940 557880 0 0 $X=301940 $Y=557500
X4431 1684 1690 111 2 1 XNR2HS $T=302560 547800 0 0 $X=302560 $Y=547420
X4432 1675 1631 1727 2 1 XNR2HS $T=306280 567960 1 0 $X=306280 $Y=562540
X4433 1705 1638 1726 2 1 XNR2HS $T=307520 557880 0 0 $X=307520 $Y=557500
X4434 1770 1592 1763 2 1 XNR2HS $T=319920 557880 0 180 $X=314340 $Y=552460
X4435 1770 1616 1790 2 1 XNR2HS $T=325500 557880 0 180 $X=319920 $Y=552460
X4436 1705 1720 1807 2 1 XNR2HS $T=327980 567960 1 180 $X=322400 $Y=567580
X4437 1705 1587 1829 2 1 XNR2HS $T=323640 567960 1 0 $X=323640 $Y=562540
X4438 1816 1611 1808 2 1 XNR2HS $T=324260 547800 0 0 $X=324260 $Y=547420
X4439 1705 1604 1851 2 1 XNR2HS $T=329220 567960 0 0 $X=329220 $Y=567580
X4440 1705 1612 1855 2 1 XNR2HS $T=329840 567960 1 0 $X=329840 $Y=562540
X4441 1816 1638 1861 2 1 XNR2HS $T=332320 557880 1 0 $X=332320 $Y=552460
X4442 1858 1631 1898 2 1 XNR2HS $T=340380 578040 1 0 $X=340380 $Y=572620
X4443 1911 1616 1892 2 1 XNR2HS $T=346580 547800 1 180 $X=341000 $Y=547420
X4444 1911 1592 1939 2 1 XNR2HS $T=345960 557880 1 0 $X=345960 $Y=552460
X4445 1905 1720 1941 2 1 XNR2HS $T=346580 567960 0 0 $X=346580 $Y=567580
X4446 1911 1611 1957 2 1 XNR2HS $T=351540 547800 0 0 $X=351540 $Y=547420
X4447 1905 1587 1981 2 1 XNR2HS $T=355880 578040 1 0 $X=355880 $Y=572620
X4448 1974 1592 1983 2 1 XNR2HS $T=356500 557880 1 0 $X=356500 $Y=552460
X4449 1974 1616 1994 2 1 XNR2HS $T=359600 547800 0 0 $X=359600 $Y=547420
X4450 1911 1638 1968 2 1 XNR2HS $T=363320 557880 1 0 $X=363320 $Y=552460
X4451 1905 1612 2023 2 1 XNR2HS $T=363940 567960 0 0 $X=363940 $Y=567580
X4452 1905 1604 2006 2 1 XNR2HS $T=363940 578040 1 0 $X=363940 $Y=572620
X4453 1945 2014 2028 2 1 XNR2HS $T=364560 608280 0 0 $X=364560 $Y=607900
X4454 1974 1611 2030 2 1 XNR2HS $T=365180 547800 0 0 $X=365180 $Y=547420
X4455 1974 1638 2043 2 1 XNR2HS $T=374480 557880 1 0 $X=374480 $Y=552460
X4456 2097 1631 2062 2 1 XNR2HS $T=381920 567960 0 180 $X=376340 $Y=562540
X4457 2065 1631 2095 2 1 XNR2HS $T=376960 567960 0 0 $X=376960 $Y=567580
X4458 2097 1587 2120 2 1 XNR2HS $T=381300 557880 0 0 $X=381300 $Y=557500
X4459 2065 1720 2109 2 1 XNR2HS $T=388120 578040 0 180 $X=382540 $Y=572620
X4460 2097 1720 2117 2 1 XNR2HS $T=385020 567960 0 0 $X=385020 $Y=567580
X4461 2065 1587 2157 2 1 XNR2HS $T=388120 578040 1 0 $X=388120 $Y=572620
X4462 2071 1604 2188 2 1 XNR2HS $T=393700 557880 0 0 $X=393700 $Y=557500
X4463 2065 1604 2204 2 1 XNR2HS $T=396180 578040 1 0 $X=396180 $Y=572620
X4464 2071 2039 2224 2 1 XNR2HS $T=399280 557880 0 0 $X=399280 $Y=557500
X4465 2321 2290 2336 2 1 XNR2HS $T=419740 557880 1 0 $X=419740 $Y=552460
X4466 2300 2327 2372 2 1 XNR2HS $T=429660 557880 1 0 $X=429660 $Y=552460
X4467 2316 2333 2406 2 1 XNR2HS $T=430900 578040 0 0 $X=430900 $Y=577660
X4468 2415 2482 2496 2 1 XNR2HS $T=447020 547800 0 0 $X=447020 $Y=547420
X4469 2641 2624 2620 2 1 XNR2HS $T=474920 648600 0 180 $X=469340 $Y=643180
X4470 2664 2651 2648 2 1 XNR2HS $T=479880 638520 1 180 $X=474300 $Y=638140
X4471 2664 2655 2654 2 1 XNR2HS $T=481120 648600 0 180 $X=475540 $Y=643180
X4472 2668 2489 2663 2 1 XNR2HS $T=482980 608280 1 180 $X=477400 $Y=607900
X4473 2664 2591 2676 2 1 XNR2HS $T=478020 658680 1 0 $X=478020 $Y=653260
X4474 2668 2546 2683 2 1 XNR2HS $T=479260 588120 0 0 $X=479260 $Y=587740
X4475 2668 2520 2686 2 1 XNR2HS $T=479880 608280 1 0 $X=479880 $Y=602860
X4476 2664 2578 2696 2 1 XNR2HS $T=481120 648600 0 0 $X=481120 $Y=648220
X4477 2668 2490 2703 2 1 XNR2HS $T=482360 618360 1 0 $X=482360 $Y=612940
X4478 2687 2517 2705 2 1 XNR2HS $T=482980 598200 0 0 $X=482980 $Y=597820
X4479 2641 2470 2710 2 1 XNR2HS $T=484220 638520 1 0 $X=484220 $Y=633100
X4480 2664 2531 2715 2 1 XNR2HS $T=484840 638520 0 0 $X=484840 $Y=638140
X4481 2664 2589 2723 2 1 XNR2HS $T=486700 648600 1 0 $X=486700 $Y=643180
X4482 2641 2521 2737 2 1 XNR2HS $T=488560 628440 1 0 $X=488560 $Y=623020
X4483 2729 2489 2749 2 1 XNR2HS $T=489800 608280 0 0 $X=489800 $Y=607900
X4484 2758 2655 2774 2 1 XNR2HS $T=493520 648600 0 0 $X=493520 $Y=648220
X4485 2687 323 2775 2 1 XNR2HS $T=494140 598200 0 0 $X=494140 $Y=597820
X4486 2729 2520 2776 2 1 XNR2HS $T=494140 608280 1 0 $X=494140 $Y=602860
X4487 2729 2490 2779 2 1 XNR2HS $T=494760 618360 1 0 $X=494760 $Y=612940
X4488 2758 2531 2780 2 1 XNR2HS $T=494760 638520 0 0 $X=494760 $Y=638140
X4489 2787 2680 2742 2 1 XNR2HS $T=500340 658680 1 180 $X=494760 $Y=658300
X4490 2787 2624 2746 2 1 XNR2HS $T=500340 668760 1 180 $X=494760 $Y=668380
X4491 2766 2521 2784 2 1 XNR2HS $T=495380 628440 1 0 $X=495380 $Y=623020
X4492 2766 2470 2785 2 1 XNR2HS $T=495380 638520 1 0 $X=495380 $Y=633100
X4493 2758 2591 2786 2 1 XNR2HS $T=495380 658680 1 0 $X=495380 $Y=653260
X4494 2766 2614 2805 2 1 XNR2HS $T=499720 608280 0 0 $X=499720 $Y=607900
X4495 2766 2589 2806 2 1 XNR2HS $T=499720 648600 1 0 $X=499720 $Y=643180
X4496 2787 2651 2781 2 1 XNR2HS $T=506540 668760 1 180 $X=500960 $Y=668380
X4497 2787 2807 2770 2 1 XNR2HS $T=507160 668760 0 180 $X=501580 $Y=663340
X4498 2766 2578 2831 2 1 XNR2HS $T=504060 658680 1 0 $X=504060 $Y=653260
X4499 2887 2490 2905 2 1 XNR2HS $T=517080 618360 1 0 $X=517080 $Y=612940
X4500 2887 2521 2923 2 1 XNR2HS $T=519560 628440 1 0 $X=519560 $Y=623020
X4501 2887 2470 2953 2 1 XNR2HS $T=525140 628440 1 0 $X=525140 $Y=623020
X4502 2887 2531 2986 2 1 XNR2HS $T=531340 628440 1 0 $X=531340 $Y=623020
X4503 3006 2589 2983 2 1 XNR2HS $T=538780 638520 1 180 $X=533200 $Y=638140
X4504 3004 2470 3023 2 1 XNR2HS $T=536920 628440 0 0 $X=536920 $Y=628060
X4505 3004 2531 3026 2 1 XNR2HS $T=538160 638520 1 0 $X=538160 $Y=633100
X4506 3006 2578 2997 2 1 XNR2HS $T=544360 648600 0 180 $X=538780 $Y=643180
X4507 3031 2624 2994 2 1 XNR2HS $T=544360 678840 0 180 $X=538780 $Y=673420
X4508 3006 3028 3042 2 1 XNR2HS $T=541260 618360 0 0 $X=541260 $Y=617980
X4509 3031 2591 3001 2 1 XNR2HS $T=546840 658680 0 180 $X=541260 $Y=653260
X4510 3038 3032 3053 2 1 XNR2HS $T=543740 578040 1 0 $X=543740 $Y=572620
X4511 3004 2589 3057 2 1 XNR2HS $T=544360 638520 1 0 $X=544360 $Y=633100
X4512 3006 2655 3021 2 1 XNR2HS $T=549940 648600 0 180 $X=544360 $Y=643180
X4513 3031 2807 3067 2 1 XNR2HS $T=553660 668760 1 180 $X=548080 $Y=668380
X4514 3031 3092 3051 2 1 XNR2HS $T=556140 678840 0 180 $X=550560 $Y=673420
X4515 3096 3032 3089 2 1 XNR2HS $T=558000 557880 1 180 $X=552420 $Y=557500
X4516 420 423 3106 2 1 XNR2HS $T=553040 547800 0 0 $X=553040 $Y=547420
X4517 3096 3092 3108 2 1 XNR2HS $T=553660 567960 1 0 $X=553660 $Y=562540
X4518 3038 3092 3076 2 1 XNR2HS $T=554280 578040 1 0 $X=554280 $Y=572620
X4519 3110 2591 3101 2 1 XNR2HS $T=559860 628440 0 180 $X=554280 $Y=623020
X4520 3031 3081 2999 2 1 XNR2HS $T=554900 668760 0 0 $X=554900 $Y=668380
X4521 3125 3081 3095 2 1 XNR2HS $T=562340 658680 0 180 $X=556760 $Y=653260
X4522 3110 2589 3123 2 1 XNR2HS $T=557380 628440 0 0 $X=557380 $Y=628060
X4523 3125 2591 3098 2 1 XNR2HS $T=563580 638520 1 180 $X=558000 $Y=638140
X4524 3125 2578 3083 2 1 XNR2HS $T=564820 638520 0 180 $X=559240 $Y=633100
X4525 3125 2655 3091 2 1 XNR2HS $T=564820 648600 0 180 $X=559240 $Y=643180
X4526 3038 3081 3136 2 1 XNR2HS $T=559860 588120 1 0 $X=559860 $Y=582700
X4527 3110 2578 3116 2 1 XNR2HS $T=560480 618360 0 0 $X=560480 $Y=617980
X4528 437 380 3077 2 1 XNR2HS $T=561720 567960 0 0 $X=561720 $Y=567580
X4529 3110 3081 3149 2 1 XNR2HS $T=563580 628440 0 0 $X=563580 $Y=628060
X4530 3156 3150 3141 2 1 XNR2HS $T=569780 638520 1 180 $X=564200 $Y=638140
X4531 3038 3150 3131 2 1 XNR2HS $T=566060 588120 1 0 $X=566060 $Y=582700
X4532 3151 3150 3167 2 1 XNR2HS $T=566680 598200 1 0 $X=566680 $Y=592780
X4533 3151 3081 3168 2 1 XNR2HS $T=566680 598200 0 0 $X=566680 $Y=597820
X4534 3151 2591 3170 2 1 XNR2HS $T=566680 608280 0 0 $X=566680 $Y=607900
X4535 3004 399 3107 2 1 XNR2HS $T=566680 618360 1 0 $X=566680 $Y=612940
X4536 3110 3150 3185 2 1 XNR2HS $T=569780 628440 0 0 $X=569780 $Y=628060
X4537 3110 2655 3099 2 1 XNR2HS $T=570400 628440 1 0 $X=570400 $Y=623020
X4538 3151 2655 3180 2 1 XNR2HS $T=573500 608280 0 0 $X=573500 $Y=607900
X4539 3156 3188 3190 2 1 XNR2HS $T=575360 648600 1 0 $X=575360 $Y=643180
X4540 3218 3092 3206 2 1 XNR2HS $T=582180 588120 1 180 $X=576600 $Y=587740
X4541 3125 3092 3163 2 1 XNR2HS $T=577220 658680 1 0 $X=577220 $Y=653260
X4542 3151 3219 3248 2 1 XNR2HS $T=582800 608280 0 0 $X=582800 $Y=607900
X4543 502 493 3242 2 1 XNR2HS $T=594580 598200 0 180 $X=589000 $Y=592780
X4544 3269 3241 3254 2 1 XNR2HS $T=594580 658680 1 180 $X=589000 $Y=658300
X4545 3207 3092 3221 2 1 XNR2HS $T=589620 628440 1 0 $X=589620 $Y=623020
X4546 3207 3188 3249 2 1 XNR2HS $T=590240 618360 0 0 $X=590240 $Y=617980
X4547 3297 3296 3280 2 1 XNR2HS $T=596440 578040 1 180 $X=590860 $Y=577660
X4548 777 4129 4122 2 1 XNR2HS $T=758260 719160 1 180 $X=752680 $Y=718780
X4549 1291 1277 1261 1 2 1252 OA12 $T=228160 699000 1 180 $X=224440 $Y=698620
X4550 46 73 1558 1 2 1568 OA12 $T=276520 578040 1 0 $X=276520 $Y=572620
X4551 1593 166 1600 1 2 172 OA12 $T=352160 578040 1 0 $X=352160 $Y=572620
X4552 211 2207 210 1 2 2248 OA12 $T=404860 578040 0 0 $X=404860 $Y=577660
X4553 292 304 305 1 2 2697 OA12 $T=481120 719160 0 0 $X=481120 $Y=718780
X4554 3442 3414 3432 1 2 3417 OA12 $T=623100 699000 0 180 $X=619380 $Y=693580
X4555 3494 3480 587 1 2 3467 OA12 $T=631780 688920 1 180 $X=628060 $Y=688540
X4556 1331 1 1333 1324 1338 1296 2 OAI22S $T=234980 699000 0 0 $X=234980 $Y=698620
X4557 24 1 1333 24 1296 1290 2 OAI22S $T=234980 709080 0 0 $X=234980 $Y=708700
X4558 24 1 1290 40 1396 43 2 OAI22S $T=246760 719160 0 0 $X=246760 $Y=718780
X4559 1430 1 1290 1430 1372 1415 2 OAI22S $T=255440 719160 0 180 $X=251720 $Y=713740
X4560 1511 1 64 62 1504 1479 2 OAI22S $T=270320 547800 1 180 $X=266600 $Y=547420
X4561 89 1 1644 96 93 78 2 OAI22S $T=295120 547800 1 180 $X=291400 $Y=547420
X4562 1645 1 1648 1653 100 1658 2 OAI22S $T=292640 557880 0 0 $X=292640 $Y=557500
X4563 92 1 99 96 98 87 2 OAI22S $T=296980 537720 1 180 $X=293260 $Y=537340
X4564 89 1 86 96 1665 1644 2 OAI22S $T=295120 547800 0 0 $X=295120 $Y=547420
X4565 1648 1 1658 1653 105 1672 2 OAI22S $T=296360 557880 0 0 $X=296360 $Y=557500
X4566 1648 1 1726 1653 1747 1727 2 OAI22S $T=310000 557880 1 0 $X=310000 $Y=552460
X4567 1729 1 1742 1733 1684 1763 2 OAI22S $T=312480 547800 0 0 $X=312480 $Y=547420
X4568 1766 1 1776 1780 1783 1771 2 OAI22S $T=315580 588120 0 0 $X=315580 $Y=587740
X4569 1795 1 1807 1761 1846 1829 2 OAI22S $T=329220 557880 0 0 $X=329220 $Y=557500
X4570 1729 1 1733 1836 1853 1742 2 OAI22S $T=330460 547800 0 0 $X=330460 $Y=547420
X4571 1795 1 1829 1761 1856 1851 2 OAI22S $T=337280 557880 1 180 $X=333560 $Y=557500
X4572 1742 1 1808 1733 1862 1861 2 OAI22S $T=334180 547800 0 0 $X=334180 $Y=547420
X4573 1835 1 1869 1543 1854 1810 2 OAI22S $T=339140 678840 1 180 $X=335420 $Y=678460
X4574 1795 1 1851 1761 149 1855 2 OAI22S $T=339760 567960 0 180 $X=336040 $Y=562540
X4575 1886 1 1861 1876 1901 1898 2 OAI22S $T=341620 567960 1 0 $X=341620 $Y=562540
X4576 1904 1 1919 1908 122 1939 2 OAI22S $T=347200 547800 0 0 $X=347200 $Y=547420
X4577 1919 1 1939 1908 163 1892 2 OAI22S $T=348440 547800 1 0 $X=348440 $Y=542380
X4578 1886 1 1898 1876 1958 1941 2 OAI22S $T=350920 567960 1 0 $X=350920 $Y=562540
X4579 1919 1 1957 1908 1962 1968 2 OAI22S $T=352160 557880 1 0 $X=352160 $Y=552460
X4580 1975 1 1941 1876 176 1981 2 OAI22S $T=357740 567960 1 0 $X=357740 $Y=562540
X4581 1973 1 2030 2043 2047 1978 2 OAI22S $T=369520 547800 1 0 $X=369520 $Y=542380
X4582 1919 1 1968 2041 190 2062 2 OAI22S $T=369520 557880 1 0 $X=369520 $Y=552460
X4583 1973 1 2043 2070 2101 2095 2 OAI22S $T=380680 557880 1 0 $X=380680 $Y=552460
X4584 2127 1 2062 2041 202 2117 2 OAI22S $T=388120 557880 0 180 $X=384400 $Y=552460
X4585 1904 1 2041 2150 2149 2127 2 OAI22S $T=388740 557880 1 0 $X=388740 $Y=552460
X4586 2100 1 2095 2109 2137 2070 2 OAI22S $T=391220 567960 1 0 $X=391220 $Y=562540
X4587 2162 1 2188 2041 2210 2224 2 OAI22S $T=400520 557880 1 0 $X=400520 $Y=552460
X4588 2100 1 2204 2070 2242 2234 2 OAI22S $T=404240 567960 0 0 $X=404240 $Y=567580
X4589 2642 1 2620 2648 2635 2605 2 OAI22S $T=473680 648600 0 0 $X=473680 $Y=648220
X4590 2642 1 2648 2654 2652 2605 2 OAI22S $T=479260 658680 1 180 $X=475540 $Y=658300
X4591 2642 1 2654 2676 2673 2605 2 OAI22S $T=483600 658680 1 180 $X=479880 $Y=658300
X4592 2688 1 2680 2620 2670 2605 2 OAI22S $T=484220 638520 1 180 $X=480500 $Y=638140
X4593 2688 1 2573 2680 2662 2605 2 OAI22S $T=485460 628440 1 180 $X=481740 $Y=628060
X4594 2583 1 2663 2686 2704 2707 2 OAI22S $T=483600 608280 0 0 $X=483600 $Y=607900
X4595 2583 1 2686 2683 2717 2712 2 OAI22S $T=486080 608280 1 0 $X=486080 $Y=602860
X4596 2583 1 2683 2705 2736 2738 2 OAI22S $T=489180 598200 0 0 $X=489180 $Y=597820
X4597 2642 1 2723 2715 2739 2713 2 OAI22S $T=489800 658680 1 0 $X=489800 $Y=653260
X4598 2583 1 2703 2663 2747 2750 2 OAI22S $T=490420 618360 1 0 $X=490420 $Y=612940
X4599 2688 1 2710 2737 2753 2713 2 OAI22S $T=491040 638520 1 0 $X=491040 $Y=633100
X4600 2688 1 2715 2710 2754 2713 2 OAI22S $T=491040 638520 0 0 $X=491040 $Y=638140
X4601 2514 1 2741 2745 2701 2762 2 OAI22S $T=491040 668760 1 0 $X=491040 $Y=663340
X4602 2734 1 2742 2746 2724 2762 2 OAI22S $T=491040 678840 1 0 $X=491040 $Y=673420
X4603 2688 1 2737 2703 2760 2713 2 OAI22S $T=492280 628440 0 0 $X=492280 $Y=628060
X4604 2741 1 2770 2742 2719 2762 2 OAI22S $T=498480 668760 0 180 $X=494760 $Y=663340
X4605 2790 1 2749 2776 2803 2775 2 OAI22S $T=500340 598200 0 0 $X=500340 $Y=597820
X4606 2790 1 2779 2749 2804 2775 2 OAI22S $T=500340 608280 1 0 $X=500340 $Y=602860
X4607 2790 1 2784 2779 2808 2775 2 OAI22S $T=501580 618360 0 0 $X=501580 $Y=617980
X4608 2790 1 2785 2784 2809 2793 2 OAI22S $T=501580 638520 1 0 $X=501580 $Y=633100
X4609 2790 1 2780 2785 2820 2793 2 OAI22S $T=503440 638520 0 0 $X=503440 $Y=638140
X4610 2741 1 2806 2780 2833 2793 2 OAI22S $T=505300 648600 1 0 $X=505300 $Y=643180
X4611 2734 1 2774 2786 2828 2762 2 OAI22S $T=505300 678840 0 0 $X=505300 $Y=678460
X4612 2741 1 2831 2806 2840 2793 2 OAI22S $T=507160 658680 0 0 $X=507160 $Y=658300
X4613 2741 1 2786 2831 2848 2793 2 OAI22S $T=508400 668760 1 0 $X=508400 $Y=663340
X4614 2932 1 2923 2905 2927 2805 2 OAI22S $T=526380 618360 0 180 $X=522660 $Y=612940
X4615 2932 1 2953 2923 2881 2805 2 OAI22S $T=530720 618360 0 180 $X=527000 $Y=612940
X4616 2932 1 2983 2986 2974 2991 2 OAI22S $T=533200 628440 0 0 $X=533200 $Y=628060
X4617 2932 1 2986 2953 2998 2991 2 OAI22S $T=533820 618360 1 0 $X=533820 $Y=612940
X4618 2981 1 2994 2999 3002 2959 2 OAI22S $T=534440 678840 1 0 $X=534440 $Y=673420
X4619 2932 1 2997 2983 2995 2991 2 OAI22S $T=538780 648600 0 180 $X=535060 $Y=643180
X4620 3010 1 3001 2997 2979 2991 2 OAI22S $T=538780 658680 0 180 $X=535060 $Y=653260
X4621 2981 1 3021 3001 2930 2959 2 OAI22S $T=542500 658680 1 180 $X=538780 $Y=658300
X4622 2981 1 2999 3021 3008 2959 2 OAI22S $T=542500 668760 0 180 $X=538780 $Y=663340
X4623 3033 1 3026 3023 3039 3042 2 OAI22S $T=543120 628440 0 0 $X=543120 $Y=628060
X4624 3025 1 2981 3037 3036 2991 2 OAI22S $T=546840 658680 1 180 $X=543120 $Y=658300
X4625 2981 1 3051 2994 3045 2959 2 OAI22S $T=548700 678840 0 180 $X=544980 $Y=673420
X4626 3033 1 3057 3026 3062 3069 2 OAI22S $T=546840 628440 0 0 $X=546840 $Y=628060
X4627 413 1 3061 3052 3063 3077 2 OAI22S $T=547460 567960 0 0 $X=547460 $Y=567580
X4628 2981 1 3067 3051 3058 2959 2 OAI22S $T=551180 668760 0 180 $X=547460 $Y=663340
X4629 3061 1 3053 3076 3080 3077 2 OAI22S $T=549320 578040 1 0 $X=549320 $Y=572620
X4630 3033 1 3083 3057 3079 3069 2 OAI22S $T=554280 638520 0 180 $X=550560 $Y=633100
X4631 3104 1 3095 3091 2992 3085 2 OAI22S $T=556140 658680 0 180 $X=552420 $Y=653260
X4632 3104 1 3091 3098 3090 3069 2 OAI22S $T=557380 648600 0 180 $X=553660 $Y=643180
X4633 3033 1 3098 3083 3056 3069 2 OAI22S $T=554900 638520 1 0 $X=554900 $Y=633100
X4634 3113 1 3089 3108 3124 3106 2 OAI22S $T=558620 557880 0 0 $X=558620 $Y=557500
X4635 3061 1 3076 3131 3133 3077 2 OAI22S $T=560480 578040 1 0 $X=560480 $Y=572620
X4636 3094 1 3116 3123 3115 3107 2 OAI22S $T=562340 618360 1 0 $X=562340 $Y=612940
X4637 3104 1 3141 3095 3138 3085 2 OAI22S $T=566680 658680 0 180 $X=562960 $Y=653260
X4638 3061 1 3131 3136 3142 3077 2 OAI22S $T=567920 578040 0 180 $X=564200 $Y=572620
X4639 458 1 3113 3130 3147 3106 2 OAI22S $T=569160 557880 0 180 $X=565440 $Y=552460
X4640 3148 1 3104 3153 3157 3085 2 OAI22S $T=566060 648600 1 0 $X=566060 $Y=643180
X4641 3104 1 3163 3141 3158 3085 2 OAI22S $T=571640 658680 0 180 $X=567920 $Y=653260
X4642 3184 1 3180 3170 3169 3172 2 OAI22S $T=574740 608280 0 180 $X=571020 $Y=602860
X4643 3104 1 3190 3163 3187 3085 2 OAI22S $T=575980 648600 1 180 $X=572260 $Y=648220
X4644 3184 1 3167 3168 3127 3172 2 OAI22S $T=572880 588120 0 0 $X=572880 $Y=587740
X4645 3184 1 3168 3180 3144 3172 2 OAI22S $T=572880 598200 1 0 $X=572880 $Y=592780
X4646 3094 1 3149 3099 3078 3186 2 OAI22S $T=572880 618360 1 0 $X=572880 $Y=612940
X4647 3094 1 3185 3149 3201 3186 2 OAI22S $T=579700 628440 1 180 $X=575980 $Y=628060
X4648 3184 1 3206 3167 3143 3172 2 OAI22S $T=580940 598200 0 180 $X=577220 $Y=592780
X4649 3094 1 3221 3185 3215 3186 2 OAI22S $T=584040 628440 1 180 $X=580320 $Y=628060
X4650 3220 1 3184 3230 3209 3242 2 OAI22S $T=581560 598200 1 0 $X=581560 $Y=592780
X4651 3184 1 3248 3206 3225 3242 2 OAI22S $T=585280 598200 0 0 $X=585280 $Y=597820
X4652 3234 1 3249 3221 3264 3186 2 OAI22S $T=585280 628440 0 0 $X=585280 $Y=628060
X4653 3192 1 3234 3268 3263 3107 2 OAI22S $T=590860 618360 0 180 $X=587140 $Y=612940
X4654 3998 1 728 4005 3020 4008 2 OAI22S $T=731600 719160 0 180 $X=727880 $Y=713740
X4655 2425 2370 2401 2 2408 2387 1 AO22 $T=437100 648600 1 0 $X=437100 $Y=643180
X4656 2470 1842 2481 2 2486 2492 1 AO22 $T=444540 628440 0 0 $X=444540 $Y=628060
X4657 2517 2216 2504 2 2469 2491 1 AO22 $T=453220 598200 1 180 $X=448260 $Y=597820
X4658 2489 2271 2500 2 2493 2512 1 AO22 $T=448260 608280 0 0 $X=448260 $Y=607900
X4659 2490 1531 2500 2 2472 2513 1 AO22 $T=448260 618360 1 0 $X=448260 $Y=612940
X4660 2520 2351 2507 2 2495 2491 1 AO22 $T=454460 608280 0 180 $X=449500 $Y=602860
X4661 2521 1576 2500 2 2505 2492 1 AO22 $T=454460 618360 1 180 $X=449500 $Y=617980
X4662 2531 1738 2481 2 2510 2492 1 AO22 $T=456320 638520 0 180 $X=451360 $Y=633100
X4663 2546 2350 2507 2 2515 2513 1 AO22 $T=458180 598200 0 180 $X=453220 $Y=592780
X4664 2591 2016 2547 2 2557 2539 1 AO22 $T=463140 618360 0 180 $X=458180 $Y=612940
X4665 2578 1840 2547 2 2558 2492 1 AO22 $T=463140 618360 1 180 $X=458180 $Y=617980
X4666 2589 1799 2481 2 2572 2492 1 AO22 $T=465620 638520 0 180 $X=460660 $Y=633100
X4667 2624 2236 2547 2 2606 2539 1 AO22 $T=471820 608280 0 180 $X=466860 $Y=602860
X4668 2651 2257 2547 2 2636 2539 1 AO22 $T=476780 608280 0 180 $X=471820 $Y=602860
X4669 2655 2081 2547 2 2634 2539 1 AO22 $T=476780 608280 1 180 $X=471820 $Y=607900
X4670 3231 2970 3243 2 3238 3265 1 AO22 $T=583420 678840 1 0 $X=583420 $Y=673420
X4671 3236 2794 3243 2 3245 3265 1 AO22 $T=584040 688920 1 0 $X=584040 $Y=683500
X4672 3165 2856 3243 2 3289 3265 1 AO22 $T=590240 688920 1 0 $X=590240 $Y=683500
X4673 3325 3241 3307 2 3240 3265 1 AO22 $T=600780 658680 1 180 $X=595820 $Y=658300
X4674 3277 2773 3243 2 3316 3265 1 AO22 $T=596440 688920 1 0 $X=596440 $Y=683500
X4675 3311 2877 3307 2 3326 3265 1 AO22 $T=598300 668760 1 0 $X=598300 $Y=663340
X4676 3315 3329 3307 2 3345 3356 1 AO22 $T=602020 618360 0 0 $X=602020 $Y=617980
X4677 3331 3064 549 2 3334 3342 1 AO22 $T=604500 638520 0 0 $X=604500 $Y=638140
X4678 3314 3369 3307 2 3366 3356 1 AO22 $T=608840 618360 0 0 $X=608840 $Y=617980
X4679 3405 3404 549 2 3400 3342 1 AO22 $T=618140 638520 0 180 $X=613180 $Y=633100
X4680 3386 3424 549 2 3410 589 1 AO22 $T=618760 608280 0 0 $X=618760 $Y=607900
X4681 3591 3601 549 2 3594 589 1 AO22 $T=649140 567960 0 0 $X=649140 $Y=567580
X4682 40 1430 1290 1409 2 1449 1 1492 MUX3 $T=257300 719160 0 0 $X=257300 $Y=718780
X4683 1648 1653 1645 1 2 104 AO12 $T=301320 557880 0 180 $X=297600 $Y=552460
X4684 1742 1733 1729 1 2 1719 AO12 $T=312480 547800 1 180 $X=308760 $Y=547420
X4685 1919 1908 1904 1 2 154 AO12 $T=347200 537720 1 180 $X=343480 $Y=537340
X4686 2669 305 314 1 2 2721 AO12 $T=485460 719160 0 0 $X=485460 $Y=718780
X4687 1772 1762 2 1787 1 1780 AOI12HS $T=316200 608280 1 0 $X=316200 $Y=602860
X4688 2397 2355 2 2369 1 2395 AOI12HS $T=432140 567960 0 180 $X=427800 $Y=562540
X4689 2415 2427 2 2447 1 2449 AOI12HS $T=438340 557880 1 0 $X=438340 $Y=552460
X4690 3269 3241 2 3239 1 3226 AOI12HS $T=587760 658680 0 180 $X=583420 $Y=653260
X4691 1469 2 61 69 1 AN2B1S $T=266600 537720 0 0 $X=266600 $Y=537340
X4692 1612 2 1795 1912 1 AN2B1S $T=342240 557880 1 0 $X=342240 $Y=552460
X4693 2039 2 1975 2048 1 AN2B1S $T=370140 567960 1 0 $X=370140 $Y=562540
X4694 2234 2 2162 2250 1 AN2B1S $T=404860 557880 1 0 $X=404860 $Y=552460
X4695 2234 2 2100 2264 1 AN2B1S $T=407960 578040 1 0 $X=407960 $Y=572620
X4696 2245 2 221 223 1 AN2B1S $T=409200 547800 0 0 $X=409200 $Y=547420
X4697 2250 2 2260 2262 1 AN2B1S $T=409200 557880 1 0 $X=409200 $Y=552460
X4698 2161 2 226 230 1 AN2B1S $T=411680 547800 1 0 $X=411680 $Y=542380
X4699 2149 2 226 2290 1 AN2B1S $T=412300 557880 1 0 $X=412300 $Y=552460
X4700 2237 2 2260 2287 1 AN2B1S $T=412300 578040 1 0 $X=412300 $Y=572620
X4701 2264 2 2260 2316 1 AN2B1S $T=417880 578040 0 0 $X=417880 $Y=577660
X4702 2573 2 2775 2684 1 AN2B1S $T=500340 628440 1 180 $X=497240 $Y=628060
X4703 2807 2 2959 2720 1 AN2B1S $T=532580 678840 0 180 $X=529480 $Y=673420
X4704 2807 2 3085 3072 1 AN2B1S $T=552420 668760 1 0 $X=552420 $Y=663340
X4705 3032 2 3077 3111 1 AN2B1S $T=555520 588120 1 0 $X=555520 $Y=582700
X4706 3032 2 3106 3129 1 AN2B1S $T=559860 567960 1 0 $X=559860 $Y=562540
X4707 3188 2 3186 3174 1 AN2B1S $T=575360 638520 1 180 $X=572260 $Y=638140
X4708 3188 2 3172 3258 1 AN2B1S $T=592720 608280 1 180 $X=589620 $Y=607900
X4709 2912 2 3426 3468 1 AN2B1S $T=629300 668760 1 0 $X=629300 $Y=663340
X4710 1404 1376 1 1282 2 1388 OAI12HS $T=251720 557880 1 180 $X=248000 $Y=557500
X4711 1490 1593 1 1600 2 1560 OAI12HS $T=282100 588120 1 0 $X=282100 $Y=582700
X4712 1535 1593 1 1600 2 1559 OAI12HS $T=283340 567960 0 0 $X=283340 $Y=567580
X4713 1592 1490 1 1616 2 1601 OAI12HS $T=286440 578040 1 0 $X=286440 $Y=572620
X4714 88 2090 1 1920 2 2130 OAI12HS $T=390600 578040 1 180 $X=386880 $Y=577660
X4715 211 210 1 1987 2 2225 OAI12HS $T=404860 578040 1 180 $X=401140 $Y=577660
X4716 2395 2393 1 2365 2 2415 OAI12HS $T=432760 557880 0 0 $X=432760 $Y=557500
X4717 2449 251 1 2439 2 257 OAI12HS $T=441440 547800 1 0 $X=441440 $Y=542380
X4718 264 266 1 2507 2 2497 OAI12HS $T=451980 567960 0 0 $X=451980 $Y=567580
X4719 3421 3469 1 3481 2 600 OAI12HS $T=627440 699000 0 0 $X=627440 $Y=698620
X4720 641 606 1 624 2 3608 OAI12HS $T=653480 537720 1 180 $X=649760 $Y=537340
X4721 18 1266 2 1290 1305 1 OR3B2S $T=228160 719160 0 0 $X=228160 $Y=718780
X4722 4421 4445 4447 2 1 835 AN3 $T=811580 567960 0 0 $X=811580 $Y=567580
X4723 4307 4455 4460 2 1 840 AN3 $T=814060 658680 0 0 $X=814060 $Y=658300
X4724 4323 4466 4470 2 1 845 AN3 $T=815920 578040 0 0 $X=815920 $Y=577660
X4725 4248 4467 4471 2 1 844 AN3 $T=815920 608280 1 0 $X=815920 $Y=602860
X4726 4190 4498 4501 2 1 855 AN3 $T=821500 608280 0 0 $X=821500 $Y=607900
X4727 4324 4504 4507 2 1 856 AN3 $T=822740 588120 0 0 $X=822740 $Y=587740
X4728 4288 4513 857 2 1 861 AN3 $T=824600 578040 1 0 $X=824600 $Y=572620
X4729 502 3192 1 2 INV3 $T=588380 578040 0 0 $X=588380 $Y=577660
X4730 3877 3855 1 2 INV3 $T=696880 598200 1 0 $X=696880 $Y=592780
X4731 1055 5406 1 2 INV3 $T=999440 658680 0 0 $X=999440 $Y=658300
X4732 5406 5358 1 2 INV3 $T=1000680 648600 0 0 $X=1000680 $Y=648220
X4733 1397 2 1401 1408 1 1414 1361 1408 1233 ICV_22 $T=249240 588120 1 0 $X=249240 $Y=582700
X4734 1421 2 1392 1428 1 1425 1451 1428 1233 ICV_22 $T=256060 648600 0 0 $X=256060 $Y=648220
X4735 1721 2 1833 1758 1 1721 1823 1712 1233 ICV_22 $T=327360 618360 1 0 $X=327360 $Y=612940
X4736 2196 2 2218 208 1 2196 2238 213 1233 ICV_22 $T=406720 688920 1 0 $X=406720 $Y=683500
X4737 2265 2 2280 229 1 2254 2291 229 1233 ICV_22 $T=412920 709080 0 0 $X=412920 $Y=708700
X4738 231 2 2417 2342 1 224 2443 233 1233 ICV_22 $T=435860 719160 1 0 $X=435860 $Y=713740
X4739 275 2 2548 277 1 2584 2574 294 1233 ICV_22 $T=462520 537720 0 0 $X=462520 $Y=537340
X4740 2436 2 2665 2725 1 2630 2752 321 1233 ICV_22 $T=489180 567960 1 0 $X=489180 $Y=562540
X4741 312 2 2812 306 1 312 2827 317 1233 ICV_22 $T=503440 557880 0 0 $X=503440 $Y=557500
X4742 2894 2 2935 360 1 2613 2961 2894 1233 ICV_22 $T=524520 578040 0 0 $X=524520 $Y=577660
X4743 406 2 496 474 1 426 3233 504 1233 ICV_22 $T=587140 537720 0 0 $X=587140 $Y=537340
X4744 3024 2 3313 3220 1 406 3296 3330 1233 ICV_22 $T=598920 588120 1 0 $X=598920 $Y=582700
X4745 3070 2 3377 3350 1 3220 3383 3148 1233 ICV_22 $T=609460 578040 1 0 $X=609460 $Y=572620
X4746 3527 2 3510 3533 1 631 3543 3480 1233 ICV_22 $T=641700 699000 1 0 $X=641700 $Y=693580
X4747 752 2 758 4049 1 759 4056 4049 1233 ICV_22 $T=739660 719160 1 0 $X=739660 $Y=713740
X4748 880 2 4583 4184 1 4184 4637 843 1233 ICV_22 $T=841960 668760 1 0 $X=841960 $Y=663340
X4749 4652 2 5498 1076 1 733 5504 1068 1233 ICV_22 $T=995720 588120 0 0 $X=995720 $Y=587740
X4750 1891 136 1818 1841 1 2 QDFFRBP $T=342240 678840 0 180 $X=329840 $Y=673420
X4751 402 385 393 331 1 2 QDFFRBP $T=543120 547800 1 0 $X=543120 $Y=542380
X4752 3463 3440 1 2 BUF2CK $T=628060 638520 0 0 $X=628060 $Y=638140
X4753 3514 3243 3505 3543 1 2 3524 AO13S $T=636740 688920 0 0 $X=636740 $Y=688540
X4754 3500 3502 2 3539 1 ND2F $T=639220 618360 0 180 $X=633020 $Y=612940
X4755 3609 3604 2 649 1 ND2F $T=655340 547800 1 180 $X=649140 $Y=547420
X4756 1348 1 1351 1278 2 ND2P $T=238700 557880 1 0 $X=238700 $Y=552460
X4757 1354 1 1346 27 2 ND2P $T=243040 537720 1 180 $X=239320 $Y=537340
X4758 1737 1 1745 1725 2 ND2P $T=310620 598200 0 0 $X=310620 $Y=597820
X4759 3216 1 3237 3272 2 ND2P $T=582800 648600 1 0 $X=582800 $Y=643180
X4760 3288 1 3272 3291 2 ND2P $T=592720 648600 0 180 $X=589000 $Y=643180
X4761 3406 1 3384 3500 2 ND2P $T=628680 618360 1 0 $X=628680 $Y=612940
X4762 3528 1 3539 3609 2 ND2P $T=652860 557880 0 180 $X=649140 $Y=552460
X4763 58 1485 1442 1 2 1478 HA1 $T=269080 668760 0 180 $X=261020 $Y=663340
X4764 1491 1481 1429 1 2 1523 HA1 $T=261640 688920 1 0 $X=261640 $Y=683500
X4765 1509 1634 1581 1 2 1586 HA1 $T=292640 688920 0 180 $X=284580 $Y=683500
X4766 1620 1628 1660 1 2 1674 HA1 $T=289540 648600 0 0 $X=289540 $Y=648220
X4767 1641 1696 1666 1 2 1663 HA1 $T=304420 628440 0 180 $X=296360 $Y=623020
X4768 1580 1740 1709 1 2 1699 HA1 $T=312480 658680 0 180 $X=304420 $Y=653260
X4769 1730 1681 1691 1 2 1714 HA1 $T=314960 618360 1 180 $X=306900 $Y=617980
X4770 1770 1773 1736 1 2 1781 HA1 $T=326120 618360 0 180 $X=318060 $Y=612940
X4771 1863 1844 1834 1 2 1830 HA1 $T=342860 608280 1 180 $X=334800 $Y=607900
X4772 1871 1913 1788 1 2 1878 HA1 $T=347200 608280 0 180 $X=339140 $Y=602860
X4773 1969 1982 1882 1 2 1954 HA1 $T=360840 598200 0 180 $X=352780 $Y=592780
X4774 2008 1988 2012 1 2 2026 HA1 $T=360220 668760 0 0 $X=360220 $Y=668380
X4775 1997 1945 2033 1 2 2015 HA1 $T=362700 598200 0 0 $X=362700 $Y=597820
X4776 2020 2012 2032 1 2 2040 HA1 $T=364560 678840 0 0 $X=364560 $Y=678460
X4777 2044 2063 1988 1 2 2031 HA1 $T=376340 668760 1 180 $X=368280 $Y=668380
X4778 2066 2033 1993 1 2 2035 HA1 $T=381300 598200 1 180 $X=373240 $Y=597820
X4779 2078 2098 2067 1 2 2061 HA1 $T=382540 658680 1 180 $X=374480 $Y=658300
X4780 2089 2067 2088 1 2 2093 HA1 $T=375720 678840 1 0 $X=375720 $Y=673420
X4781 2101 1853 2103 1 2 2122 HA1 $T=378200 547800 0 0 $X=378200 $Y=547420
X4782 2108 2088 2063 1 2 2124 HA1 $T=378820 668760 0 0 $X=378820 $Y=668380
X4783 2164 2183 2098 1 2 2142 HA1 $T=397420 668760 0 180 $X=389360 $Y=663340
X4784 2166 2184 2152 1 2 205 HA1 $T=397420 719160 0 180 $X=389360 $Y=713740
X4785 2177 2154 2183 1 2 2198 HA1 $T=390600 668760 0 0 $X=390600 $Y=668380
X4786 2218 2235 2199 1 2 2197 HA1 $T=406720 699000 1 180 $X=398660 $Y=698620
X4787 2222 2238 2205 1 2 2203 HA1 $T=407340 678840 1 180 $X=399280 $Y=678460
X4788 2192 2210 2245 1 2 2247 HA1 $T=400520 547800 0 0 $X=400520 $Y=547420
X4789 2209 2217 2244 1 2 2255 HA1 $T=401140 658680 1 0 $X=401140 $Y=653260
X4790 2231 2241 2214 1 2 2213 HA1 $T=409200 709080 1 180 $X=401140 $Y=708700
X4791 2221 2258 2217 1 2 2226 HA1 $T=411060 658680 1 180 $X=403000 $Y=658300
X4792 2246 2249 6233 1 2 2211 HA1 $T=413540 678840 0 180 $X=405480 $Y=673420
X4793 2268 2244 2285 1 2 2306 HA1 $T=408580 648600 0 0 $X=408580 $Y=648220
X4794 2269 2275 2258 1 2 2330 HA1 $T=412300 658680 1 0 $X=412300 $Y=653260
X4795 2288 2310 2275 1 2 2273 HA1 $T=420360 668760 0 180 $X=412300 $Y=663340
X4796 2295 2279 2311 1 2 2324 HA1 $T=412920 678840 0 0 $X=412920 $Y=678460
X4797 2296 2276 2297 1 2 2326 HA1 $T=413540 699000 1 0 $X=413540 $Y=693580
X4798 2303 2278 2319 1 2 2331 HA1 $T=414160 567960 0 0 $X=414160 $Y=567580
X4799 2291 2289 2323 1 2 235 HA1 $T=414780 719160 1 0 $X=414780 $Y=713740
X4800 2280 2293 2339 1 2 2348 HA1 $T=416640 709080 0 0 $X=416640 $Y=708700
X4801 2329 2353 2310 1 2 2314 HA1 $T=427180 648600 0 180 $X=419120 $Y=643180
X4802 2335 2320 2354 1 2 2367 HA1 $T=419740 668760 0 0 $X=419740 $Y=668380
X4803 2396 2346 2353 1 2 2408 HA1 $T=427180 638520 0 0 $X=427180 $Y=638140
X4804 2373 2285 2407 1 2 2402 HA1 $T=428420 648600 0 0 $X=428420 $Y=648220
X4805 2419 2409 2446 1 2 2486 HA1 $T=434620 638520 1 0 $X=434620 $Y=633100
X4806 2418 2421 2441 1 2 2472 HA1 $T=436480 618360 0 0 $X=436480 $Y=617980
X4807 2432 2407 2454 1 2 2442 HA1 $T=436480 658680 1 0 $X=436480 $Y=653260
X4808 2444 2426 6234 1 2 2469 HA1 $T=437100 598200 0 0 $X=437100 $Y=597820
X4809 2466 2445 2465 1 2 2495 HA1 $T=439580 608280 1 0 $X=439580 $Y=602860
X4810 2428 2441 2445 1 2 2493 HA1 $T=439580 618360 1 0 $X=439580 $Y=612940
X4811 2473 2446 2421 1 2 2505 HA1 $T=440820 628440 1 0 $X=440820 $Y=623020
X4812 2435 2450 6235 1 2 2484 HA1 $T=440820 638520 0 0 $X=440820 $Y=638140
X4813 2483 2465 2426 1 2 2515 HA1 $T=442680 598200 1 0 $X=442680 $Y=592780
X4814 2508 2454 2519 1 2 2487 HA1 $T=447640 658680 1 0 $X=447640 $Y=653260
X4815 2506 2556 2409 1 2 2510 HA1 $T=460040 628440 1 180 $X=451980 $Y=628060
X4816 2540 2564 2450 1 2 2518 HA1 $T=461900 638520 1 180 $X=453840 $Y=638140
X4817 2541 2519 2564 1 2 2561 HA1 $T=454460 648600 0 0 $X=454460 $Y=648220
X4818 2530 2431 2575 1 2 2586 HA1 $T=456320 598200 0 0 $X=456320 $Y=597820
X4819 2560 2607 2576 1 2 2557 HA1 $T=469340 608280 1 180 $X=461280 $Y=607900
X4820 2587 2609 2556 1 2 2572 HA1 $T=469340 628440 1 180 $X=461280 $Y=628060
X4821 2535 2576 2609 1 2 2558 HA1 $T=464380 618360 0 0 $X=464380 $Y=617980
X4822 2598 2585 2579 1 2 2455 HA1 $T=472440 658680 0 180 $X=464380 $Y=653260
X4823 2599 2575 2623 1 2 2606 HA1 $T=465000 598200 0 0 $X=465000 $Y=597820
X4824 2610 2603 6236 1 2 2590 HA1 $T=473060 638520 1 180 $X=465000 $Y=638140
X4825 2644 2662 2625 1 2 6237 HA1 $T=479260 628440 1 180 $X=471200 $Y=628060
X4826 2622 2647 2607 1 2 2634 HA1 $T=480500 618360 0 180 $X=472440 $Y=612940
X4827 2660 2623 2647 1 2 2636 HA1 $T=482360 598200 1 180 $X=474300 $Y=597820
X4828 2701 2719 2685 1 2 2677 HA1 $T=490420 668760 0 180 $X=482360 $Y=663340
X4829 3036 3058 3027 1 2 2763 HA1 $T=549320 678840 1 180 $X=541260 $Y=678460
X4830 3063 3080 3049 1 2 3044 HA1 $T=553660 588120 0 180 $X=545600 $Y=582700
X4831 3152 3139 3162 1 2 467 HA1 $T=563580 547800 0 0 $X=563580 $Y=547420
X4832 3147 3124 6238 1 2 3173 HA1 $T=563580 557880 0 0 $X=563580 $Y=557500
X4833 3157 3187 3164 1 2 3022 HA1 $T=578460 658680 1 180 $X=570400 $Y=658300
X4834 3209 3225 3118 1 2 3200 HA1 $T=584040 598200 1 180 $X=575980 $Y=597820
X4835 3191 3199 3223 1 2 3235 HA1 $T=576600 578040 1 0 $X=576600 $Y=572620
X4836 3196 3233 481 1 2 478 HA1 $T=585280 537720 1 180 $X=577220 $Y=537340
X4837 3263 3264 3256 1 2 3160 HA1 $T=596440 638520 0 180 $X=588380 $Y=633100
X4838 1491 1509 1518 2 1 XOR2HS $T=267220 557880 1 0 $X=267220 $Y=552460
X4839 1578 1509 1552 2 1 XOR2HS $T=282100 547800 1 180 $X=276520 $Y=547420
X4840 1578 1580 1633 2 1 XOR2HS $T=287680 567960 0 0 $X=287680 $Y=567580
X4841 1641 1580 1659 2 1 XOR2HS $T=292020 578040 1 0 $X=292020 $Y=572620
X4842 1641 1730 1744 2 1 XOR2HS $T=308760 567960 0 0 $X=308760 $Y=567580
X4843 1770 1730 1786 2 1 XOR2HS $T=315580 567960 0 0 $X=315580 $Y=567580
X4844 1858 1863 1877 2 1 XOR2HS $T=336040 578040 0 0 $X=336040 $Y=577660
X4845 1871 1863 1937 2 1 XOR2HS $T=345340 578040 0 0 $X=345340 $Y=577660
X4846 1871 1969 1977 2 1 XOR2HS $T=354640 578040 0 0 $X=354640 $Y=577660
X4847 2066 1969 2049 2 1 XOR2HS $T=378200 578040 0 180 $X=372620 $Y=572620
X4848 2400 2375 2416 2 1 XOR2HS $T=432760 567960 0 0 $X=432760 $Y=567580
X4849 2395 2412 2440 2 1 XOR2HS $T=436480 567960 1 0 $X=436480 $Y=562540
X4850 2449 2438 255 2 1 XOR2HS $T=440820 537720 0 0 $X=440820 $Y=537340
X4851 2525 2523 263 2 1 XOR2HS $T=456320 547800 0 180 $X=450740 $Y=542380
X4852 2524 2526 2538 2 1 XOR2HS $T=453840 557880 0 0 $X=453840 $Y=557500
X4853 2538 2545 270 2 1 XOR2HS $T=456320 567960 1 0 $X=456320 $Y=562540
X4854 2566 2562 2543 2 1 XOR2HS $T=461900 578040 1 180 $X=456320 $Y=577660
X4855 2571 2543 2545 2 1 XOR2HS $T=462520 578040 0 180 $X=456940 $Y=572620
X4856 2574 2570 2553 2 1 XOR2HS $T=463140 547800 0 180 $X=457560 $Y=542380
X4857 2632 2596 285 2 1 XOR2HS $T=473680 547800 1 180 $X=468100 $Y=547420
X4858 2638 2592 286 2 1 XOR2HS $T=474300 547800 0 180 $X=468720 $Y=542380
X4859 2643 2639 2526 2 1 XOR2HS $T=475540 557880 1 180 $X=469960 $Y=557500
X4860 2621 2649 2661 2 1 XOR2HS $T=474300 588120 1 0 $X=474300 $Y=582700
X4861 2667 2665 2571 2 1 XOR2HS $T=481120 578040 0 180 $X=475540 $Y=572620
X4862 2640 2661 307 2 1 XOR2HS $T=480500 588120 1 0 $X=480500 $Y=582700
X4863 2702 2699 2666 2 1 XOR2HS $T=487320 578040 0 180 $X=481740 $Y=572620
X4864 2692 2726 2744 2 1 XOR2HS $T=489180 567960 0 0 $X=489180 $Y=567580
X4865 2752 2718 2726 2 1 XOR2HS $T=492900 557880 0 0 $X=492900 $Y=557500
X4866 2800 2797 2783 2 1 XOR2HS $T=503440 578040 1 180 $X=497860 $Y=577660
X4867 2783 2791 336 2 1 XOR2HS $T=499100 578040 1 0 $X=499100 $Y=572620
X4868 2744 2799 2810 2 1 XOR2HS $T=500960 567960 1 0 $X=500960 $Y=562540
X4869 2768 2801 2814 2 1 XOR2HS $T=501580 547800 0 0 $X=501580 $Y=547420
X4870 2729 323 2825 2 1 XOR2HS $T=503440 598200 1 0 $X=503440 $Y=592780
X4871 2814 2843 2857 2 1 XOR2HS $T=509640 557880 1 0 $X=509640 $Y=552460
X4872 2846 2835 2801 2 1 XOR2HS $T=510260 547800 1 0 $X=510260 $Y=542380
X4873 2865 2863 2849 2 1 XOR2HS $T=515840 567960 0 180 $X=510260 $Y=562540
X4874 2849 2829 2870 2 1 XOR2HS $T=511500 557880 0 0 $X=511500 $Y=557500
X4875 2966 2960 2951 2 1 XOR2HS $T=533200 567960 1 180 $X=527620 $Y=567580
X4876 2870 2941 2964 2 1 XOR2HS $T=528240 557880 0 0 $X=528240 $Y=557500
X4877 2951 2857 2972 2 1 XOR2HS $T=529480 557880 1 0 $X=529480 $Y=552460
X4878 2812 2943 2996 2 1 XOR2HS $T=532580 567960 1 0 $X=532580 $Y=562540
X4879 3009 2996 2985 2 1 XOR2HS $T=539400 567960 1 180 $X=533820 $Y=567580
X4880 2646 346 2967 2 1 XOR2HS $T=540640 588120 0 180 $X=535060 $Y=582700
X4881 2985 2810 2989 2 1 XOR2HS $T=538780 567960 1 0 $X=538780 $Y=562540
X4882 3004 3028 3073 2 1 XOR2HS $T=547460 618360 0 0 $X=547460 $Y=617980
X4883 420 380 3103 2 1 XOR2HS $T=552420 567960 0 0 $X=552420 $Y=567580
X4884 3096 423 3122 2 1 XOR2HS $T=557380 547800 1 0 $X=557380 $Y=542380
X4885 3207 399 3217 2 1 XOR2HS $T=577220 618360 1 0 $X=577220 $Y=612940
X4886 3218 493 3262 2 1 XOR2HS $T=584660 588120 1 0 $X=584660 $Y=582700
X4887 1549 1608 1590 1 2 1534 MAO222 $T=288920 648600 1 180 $X=283960 $Y=648220
X4888 1607 1614 1583 1 2 1599 MAO222 $T=289540 608280 0 180 $X=284580 $Y=602860
X4889 1618 1619 1599 1 2 1590 MAO222 $T=286440 638520 1 0 $X=286440 $Y=633100
X4890 1622 1646 1655 1 2 1583 MAO222 $T=295740 608280 0 180 $X=290780 $Y=602860
X4891 1654 52 1664 1 2 1668 MAO222 $T=293260 699000 1 0 $X=293260 $Y=693580
X4892 1635 1501 1685 1 2 1664 MAO222 $T=301320 688920 1 180 $X=296360 $Y=688540
X4893 1657 1500 1668 1 2 1688 MAO222 $T=296980 709080 0 0 $X=296980 $Y=708700
X4894 1697 108 1688 1 2 112 MAO222 $T=301320 719160 0 0 $X=301320 $Y=718780
X4895 1706 55 1713 1 2 1685 MAO222 $T=306900 688920 0 180 $X=301940 $Y=683500
X4896 1669 1683 1725 1 2 1655 MAO222 $T=310000 598200 1 180 $X=305040 $Y=597820
X4897 56 109 119 1 2 128 MAO222 $T=311240 719160 1 0 $X=311240 $Y=713740
X4898 1765 1760 1703 1 2 1713 MAO222 $T=317440 688920 0 180 $X=312480 $Y=683500
X4899 1784 1788 1791 1 2 1766 MAO222 $T=316820 598200 1 0 $X=316820 $Y=592780
X4900 1681 1806 1811 1 2 1822 MAO222 $T=320540 688920 0 0 $X=320540 $Y=688540
X4901 1930 1935 1948 1 2 1923 MAO222 $T=352160 688920 0 180 $X=347200 $Y=683500
X4902 1985 1925 1982 1 2 1964 MAO222 $T=365180 618360 1 180 $X=360220 $Y=617980
X4903 3371 3403 3415 1 2 3448 MAO222 $T=620000 578040 1 0 $X=620000 $Y=572620
X4904 1313 1289 1246 2 1 1237 XOR3 $T=231260 578040 0 180 $X=220100 $Y=572620
X4905 1299 1274 1248 2 1 1234 XOR3 $T=231260 668760 0 180 $X=220100 $Y=663340
X4906 1308 1292 1255 2 1 1241 XOR3 $T=231880 628440 1 180 $X=220720 $Y=628060
X4907 1311 1293 1256 2 1 1236 XOR3 $T=231880 668760 1 180 $X=220720 $Y=668380
X4908 1309 1294 1257 2 1 1242 XOR3 $T=231880 678840 0 180 $X=220720 $Y=673420
X4909 1269 1273 1315 2 1 1319 XOR3 $T=223820 608280 0 0 $X=223820 $Y=607900
X4910 1317 1318 1278 2 1 1267 XOR3 $T=236220 547800 1 180 $X=225060 $Y=547420
X4911 1344 1349 1304 2 1 1295 XOR3 $T=241180 618360 0 180 $X=230020 $Y=612940
X4912 1336 1352 1323 2 1 1314 XOR3 $T=244900 567960 1 180 $X=233740 $Y=567580
X4913 1325 1322 1337 2 1 1302 XOR3 $T=248000 598200 0 180 $X=236840 $Y=592780
X4914 1522 1527 1512 2 1 1502 XOR3 $T=279000 658680 1 180 $X=267840 $Y=658300
X4915 1526 1521 1534 2 1 1525 XOR3 $T=282720 648600 1 180 $X=271560 $Y=648220
X4916 1607 1614 1583 2 1 1572 XOR3 $T=291400 598200 1 180 $X=280240 $Y=597820
X4917 1549 1608 1590 2 1 1574 XOR3 $T=292640 638520 1 180 $X=281480 $Y=638140
X4918 1618 1619 1599 2 1 1577 XOR3 $T=295120 628440 0 180 $X=283960 $Y=623020
X4919 1622 1646 1655 2 1 1642 XOR3 $T=292640 598200 0 0 $X=292640 $Y=597820
X4920 1669 1683 1725 2 1 1734 XOR3 $T=299460 598200 1 0 $X=299460 $Y=592780
X4921 1784 1788 1791 2 1 1866 XOR3 $T=322400 598200 1 0 $X=322400 $Y=592780
X4922 1681 1806 1811 2 1 146 XOR3 $T=322400 699000 1 0 $X=322400 $Y=693580
X4923 1930 1935 1948 2 1 180 XOR3 $T=352160 688920 1 0 $X=352160 $Y=683500
X4924 2970 3189 3177 2 1 3238 XOR3 $T=572880 668760 0 0 $X=572880 $Y=668380
X4925 2830 3229 3228 2 1 3289 XOR3 $T=587140 699000 0 0 $X=587140 $Y=698620
X4926 2877 3250 3260 2 1 3326 XOR3 $T=590240 668760 0 0 $X=590240 $Y=668380
X4927 3064 3283 3291 2 1 3334 XOR3 $T=591480 638520 0 0 $X=591480 $Y=638140
X4928 2773 3261 3251 2 1 3316 XOR3 $T=591480 688920 0 0 $X=591480 $Y=688540
X4929 3303 3306 3339 2 1 3345 XOR3 $T=597060 628440 1 0 $X=597060 $Y=623020
X4930 3369 3412 3379 2 1 3366 XOR3 $T=620620 628440 0 180 $X=609460 $Y=623020
X4931 3371 3403 3415 2 1 3446 XOR3 $T=615660 567960 1 0 $X=615660 $Y=562540
X4932 3440 3438 3320 2 1 3400 XOR3 $T=628060 638520 1 180 $X=616900 $Y=638140
X4933 3406 3444 3384 2 1 3410 XOR3 $T=628680 618360 1 180 $X=617520 $Y=617980
X4934 3528 3531 3539 2 1 3594 XOR3 $T=636740 567960 0 0 $X=636740 $Y=567580
X4935 1669 1714 2 1724 1679 1 1646 FA1 $T=297600 608280 1 0 $X=297600 $Y=602860
X4936 1772 1823 2 1834 1781 1 1683 FA1 $T=316200 608280 0 0 $X=316200 $Y=607900
X4937 155 1740 2 1785 1822 1 1748 FA1 $T=343480 688920 1 180 $X=327980 $Y=688540
X4938 1942 1878 2 1882 1932 1 1791 FA1 $T=350300 598200 1 180 $X=334800 $Y=597820
X4939 161 1844 2 1873 1923 1 1811 FA1 $T=350300 699000 0 180 $X=334800 $Y=693580
X4940 1970 1954 2 1928 1993 1 1932 FA1 $T=363940 608280 0 180 $X=348440 $Y=602860
X4941 348 2895 2 2904 2860 1 6239 FA1 $T=509020 608280 1 0 $X=509020 $Y=602860
X4942 505 3253 2 3308 527 1 3348 FA1 $T=590860 537720 0 0 $X=590860 $Y=537340
X4943 3355 3213 2 3279 3287 1 3278 FA1 $T=606360 567960 0 180 $X=590860 $Y=562540
X4944 3401 3335 2 3328 3338 1 3304 FA1 $T=613800 557880 1 180 $X=598300 $Y=557500
X4945 568 3355 2 3391 3348 1 604 FA1 $T=613800 537720 0 0 $X=613800 $Y=537340
X4946 3391 3270 2 3445 3401 1 3490 FA1 $T=616280 557880 0 0 $X=616280 $Y=557500
X4947 3519 3305 2 3385 3425 1 3419 FA1 $T=634260 578040 1 180 $X=618760 $Y=577660
X4948 606 3474 2 3525 609 1 638 FA1 $T=631780 537720 0 0 $X=631780 $Y=537340
X4949 610 3278 2 3490 3580 1 637 FA1 $T=633020 547800 0 0 $X=633020 $Y=547420
X4950 624 3538 2 3563 3535 1 641 FA1 $T=639840 547800 1 0 $X=639840 $Y=542380
X4951 3011 2875 2 1 2969 390 2889 2962 397 3016 2984 1233 ICV_24 $T=538780 709080 1 180 $X=534440 $Y=708700
X4952 3849 3856 2 1 3800 3826 3855 3859 3813 3861 3482 1233 ICV_24 $T=695020 588120 1 180 $X=690680 $Y=587740
X4953 3975 3856 2 1 3947 715 3855 3903 3983 3976 3930 1233 ICV_24 $T=722300 567960 1 180 $X=717960 $Y=567580
X4954 4228 4153 2 1 4205 663 4148 4168 4211 4193 4227 1233 ICV_24 $T=770040 638520 0 180 $X=765700 $Y=633100
X4955 4273 4020 2 1 4239 4253 4258 4254 4182 4274 4242 1233 ICV_24 $T=779340 608280 1 180 $X=775000 $Y=607900
X4956 4330 4153 2 1 4329 4326 4283 4294 4350 4353 4305 1233 ICV_24 $T=792980 648600 0 180 $X=788640 $Y=643180
X4957 4358 4153 2 1 4308 4068 4283 4294 4322 4373 4367 1233 ICV_24 $T=796080 648600 1 180 $X=791740 $Y=648220
X4958 4580 4528 2 1 4552 4557 4566 4561 4589 4535 4572 1233 ICV_24 $T=835760 678840 0 180 $X=831420 $Y=673420
X4959 4702 897 2 1 4669 4537 4708 4718 4642 4724 903 1233 ICV_24 $T=856220 598200 1 180 $X=851880 $Y=597820
X4960 4706 891 2 1 4675 4625 892 901 4647 4730 4676 1233 ICV_24 $T=856840 547800 1 180 $X=852500 $Y=547420
X4961 4984 4989 2 1 4948 821 4963 4573 4991 4962 5010 1233 ICV_24 $T=905200 668760 0 180 $X=900860 $Y=663340
X4962 5050 4925 2 1 5031 965 4912 4786 5043 5040 5060 1233 ICV_24 $T=915120 598200 1 180 $X=910780 $Y=597820
X4963 5471 5408 2 1 5475 5458 5424 5403 5511 5438 1080 1233 ICV_24 $T=998820 588120 0 180 $X=994480 $Y=582700
X4964 5488 5608 2 1 5731 5732 5512 5755 5741 5759 5766 1233 ICV_24 $T=1040980 628440 1 180 $X=1036640 $Y=628060
X4965 5877 5806 2 1 5841 5858 5829 5554 5880 5866 5894 1233 ICV_24 $T=1063920 699000 0 180 $X=1059580 $Y=693580
X4966 5956 5887 2 1 5924 5890 5693 5911 5899 5957 5909 1233 ICV_24 $T=1079420 668760 0 180 $X=1075080 $Y=663340
X4967 6111 5751 2 1 6072 6056 5868 5861 6014 6091 6125 1233 ICV_24 $T=1107320 588120 0 180 $X=1102980 $Y=582700
X4968 1917 1 2 2148 2216 2148 2167 22 1233 ICV_25 $T=395560 608280 0 0 $X=395560 $Y=607900
X4969 2208 1 2 2298 2351 2298 2292 20 1233 ICV_25 $T=418500 608280 0 0 $X=418500 $Y=607900
X4970 3284 1 2 676 3504 3587 3761 678 1233 ICV_25 $T=678900 709080 0 0 $X=678900 $Y=708700
X4971 3824 1 2 4037 4078 4048 4057 655 1233 ICV_25 $T=735320 668760 0 0 $X=735320 $Y=668380
X4972 4116 1 2 767 4143 4075 4100 767 1233 ICV_25 $T=748340 588120 0 0 $X=748340 $Y=587740
X4973 4168 1 2 4294 4317 4104 4262 4253 1233 ICV_25 $T=780580 648600 1 0 $X=780580 $Y=643180
X4974 4169 1 2 938 4946 899 939 936 1233 ICV_25 $T=890320 719160 0 0 $X=890320 $Y=718780
X4975 4767 1 2 4969 4993 4925 4968 4969 1233 ICV_25 $T=899620 618360 0 0 $X=899620 $Y=617980
X4976 4515 1 2 5131 5183 4955 5146 5131 1233 ICV_25 $T=936200 628440 1 0 $X=936200 $Y=623020
X4977 5381 1 2 5396 5429 5412 5335 816 1233 ICV_25 $T=979600 628440 0 0 $X=979600 $Y=628060
X4978 5445 1 2 5458 5485 5345 5411 5458 1233 ICV_25 $T=988900 588120 0 0 $X=988900 $Y=587740
X4979 5742 1 2 5750 5761 5605 5708 1118 1233 ICV_25 $T=1039120 709080 0 0 $X=1039120 $Y=708700
X4980 5578 1 2 5853 5852 5853 5836 5858 1233 ICV_25 $T=1057100 678840 0 0 $X=1057100 $Y=678460
X4981 5579 1 2 5887 5912 5812 5889 5890 1233 ICV_25 $T=1063300 668760 1 0 $X=1063300 $Y=663340
X4982 1140 1 2 5910 5945 5782 5928 5910 1233 ICV_25 $T=1070740 598200 1 0 $X=1070740 $Y=592780
X4983 5932 1 2 6002 6017 5782 5976 6005 1233 ICV_25 $T=1086860 588120 0 0 $X=1086860 $Y=587740
X4984 1143 1 2 1160 1168 5842 6028 1164 1233 ICV_25 $T=1091200 547800 1 0 $X=1091200 $Y=542380
X4985 1824 1536 2 1 1803 1620 1799 1536 1782 1641 1233 ICV_26 $T=322400 618360 1 180 $X=318060 $Y=617980
X4986 2219 2163 2 1 2111 159 2182 2163 2151 1587 1233 ICV_26 $T=396800 638520 0 180 $X=392460 $Y=633100
X4987 2334 2298 2 1 2313 2014 2305 2298 2284 165 1233 ICV_26 $T=419120 628440 0 180 $X=414780 $Y=623020
X4988 2864 2875 2 1 2735 343 2817 2839 2796 340 1233 ICV_26 $T=510260 709080 1 180 $X=505920 $Y=708700
X4989 3949 3776 2 1 3961 715 3959 3792 3923 715 1233 ICV_26 $T=719200 588120 1 180 $X=714860 $Y=587740
X4990 4149 4037 2 1 4102 4107 4124 4048 4097 4107 1233 ICV_26 $T=750820 668760 1 180 $X=746480 $Y=668380
X4991 4209 4095 2 1 4165 4183 4181 4043 4096 4116 1233 ICV_26 $T=760740 598200 1 180 $X=756400 $Y=597820
X4992 3312 4108 2 1 4235 4210 3416 4108 4219 796 1233 ICV_26 $T=777480 678840 0 180 $X=773140 $Y=673420
X4993 3372 4066 2 1 4389 819 4387 4066 4315 796 1233 ICV_26 $T=802900 709080 1 180 $X=798560 $Y=708700
X4994 4574 4530 2 1 4485 4525 4554 4487 4484 4525 1233 ICV_26 $T=830800 588120 1 180 $X=826460 $Y=587740
X4995 4712 897 2 1 4666 4525 4682 891 4655 4525 1233 ICV_26 $T=853120 588120 1 180 $X=848780 $Y=587740
X4996 905 899 2 1 902 819 4723 899 4684 871 1233 ICV_26 $T=858080 719160 1 180 $X=853740 $Y=718780
X4997 4776 913 2 1 4754 4674 909 891 4681 4674 1233 ICV_26 $T=864280 598200 1 180 $X=859940 $Y=597820
X4998 5828 5578 2 1 5803 5781 5800 5590 5780 5781 1233 ICV_26 $T=1050280 678840 1 180 $X=1045940 $Y=678460
X4999 5963 5838 2 1 5923 5946 5898 5838 5882 5897 1233 ICV_26 $T=1076940 628440 1 180 $X=1072600 $Y=628060
X5000 5992 5845 2 1 5944 5650 5970 5853 5883 5650 1233 ICV_26 $T=1083140 648600 1 180 $X=1078800 $Y=648220
X5001 4745 2 1 910 BUF3 $T=864900 628440 0 0 $X=864900 $Y=628060
X5002 5358 2 1 1039 BUF3 $T=980840 567960 0 0 $X=980840 $Y=567580
X5003 3481 3421 3503 1 2 1916 AN3S $T=635500 699000 1 180 $X=631780 $Y=698620
X5004 4403 4433 4434 1 2 829 AN3S $T=809100 678840 1 0 $X=809100 $Y=673420
X5005 4430 4438 4440 1 2 831 AN3S $T=810340 658680 0 0 $X=810340 $Y=658300
X5006 4359 4451 4452 1 2 838 AN3S $T=812820 668760 0 0 $X=812820 $Y=668380
X5007 4017 4490 4493 1 2 850 AN3S $T=819640 668760 0 0 $X=819640 $Y=668380
X5008 4009 4526 4531 1 2 864 AN3S $T=825840 608280 0 0 $X=825840 $Y=607900
X5009 4406 4437 2 4398 4441 1 OR3B2 $T=809100 678840 0 0 $X=809100 $Y=678460
X5010 3855 1 699 2 BUF4CK $T=704320 557880 1 0 $X=704320 $Y=552460
X5011 1629 1849 1896 1899 2 1906 1 AOI13HS $T=342240 678840 0 0 $X=342240 $Y=678460
X5012 3494 3578 636 3510 2 3543 1 AOI13HS $T=647280 688920 1 180 $X=643560 $Y=688540
X5013 3528 3531 2 3539 3604 3531 1 AOI22HT $T=636740 567960 1 0 $X=636740 $Y=562540
X5014 1274 1299 1248 1255 1 2 MAO222P $T=230020 658680 0 0 $X=230020 $Y=658300
X5015 1322 1325 1337 1246 1 2 MAO222P $T=237460 588120 1 180 $X=231880 $Y=587740
X5016 1292 1308 1255 1304 1 2 MAO222P $T=232500 638520 1 0 $X=232500 $Y=633100
X5017 1293 1311 1256 1248 1 2 MAO222P $T=233120 668760 0 0 $X=233120 $Y=668380
X5018 1289 1313 1246 1323 1 2 MAO222P $T=233740 578040 1 0 $X=233740 $Y=572620
X5019 1294 1309 1257 1256 1 2 MAO222P $T=240560 678840 0 180 $X=234980 $Y=673420
X5020 1273 1269 1315 1337 1 2 MAO222P $T=243660 608280 0 180 $X=238080 $Y=602860
X5021 1349 1344 1304 1315 1 2 MAO222P $T=242420 618360 1 0 $X=242420 $Y=612940
X5022 1521 1526 1534 1512 1 2 MAO222P $T=274040 658680 0 180 $X=268460 $Y=653260
X5023 1527 1522 1512 1257 1 2 MAO222P $T=270320 668760 1 0 $X=270320 $Y=663340
X5024 3229 2830 3228 3251 1 2 MAO222P $T=581560 699000 0 0 $X=581560 $Y=698620
X5025 3250 2851 3260 3177 1 2 MAO222P $T=584660 668760 0 0 $X=584660 $Y=668380
X5026 3261 2773 3251 3260 1 2 MAO222P $T=585900 688920 0 0 $X=585900 $Y=688540
X5027 3283 3064 3291 3320 1 2 MAO222P $T=593960 648600 1 0 $X=593960 $Y=643180
X5028 3412 3369 3379 3339 1 2 MAO222P $T=620620 628440 1 180 $X=615040 $Y=628060
X5029 3438 3440 3320 3379 1 2 MAO222P $T=624960 638520 0 180 $X=619380 $Y=633100
X5030 1329 1 2 1307 1265 1286 1233 ICV_27 $T=237460 588120 0 0 $X=237460 $Y=587740
X5031 1657 1 2 1662 1635 1682 1233 ICV_27 $T=295120 709080 1 0 $X=295120 $Y=703660
X5032 1703 1 2 1723 1706 1751 1233 ICV_27 $T=306900 678840 1 0 $X=306900 $Y=673420
X5033 1842 1 2 1824 1825 1848 1233 ICV_27 $T=331080 618360 0 0 $X=331080 $Y=617980
X5034 2058 1 2 2059 2082 2073 1233 ICV_27 $T=373240 618360 0 0 $X=373240 $Y=617980
X5035 2091 1 2 2110 2106 2118 1233 ICV_27 $T=379440 588120 0 0 $X=379440 $Y=587740
X5036 2111 1 2 2136 2107 2145 1233 ICV_27 $T=383780 618360 0 0 $X=383780 $Y=617980
X5037 2767 1 2 2794 2798 2821 1233 ICV_27 $T=496620 678840 1 0 $X=496620 $Y=673420
X5038 335 1 2 342 345 354 1233 ICV_27 $T=502200 688920 0 0 $X=502200 $Y=688540
X5039 357 1 2 365 2885 2914 1233 ICV_27 $T=512120 678840 0 0 $X=512120 $Y=678460
X5040 381 1 2 387 388 394 1233 ICV_27 $T=528240 668760 0 0 $X=528240 $Y=668380
X5041 3018 1 2 3035 3041 3068 1233 ICV_27 $T=539400 648600 0 0 $X=539400 $Y=648220
X5042 439 1 2 449 457 468 1233 ICV_27 $T=562960 588120 0 0 $X=562960 $Y=587740
X5043 3204 1 2 3255 503 511 1233 ICV_27 $T=584660 699000 1 0 $X=584660 $Y=693580
X5044 3286 1 2 3302 522 536 1233 ICV_27 $T=592720 598200 0 0 $X=592720 $Y=597820
X5045 533 1 2 545 551 561 1233 ICV_27 $T=601400 608280 0 0 $X=601400 $Y=607900
X5046 547 1 2 560 562 576 1233 ICV_27 $T=605740 648600 0 0 $X=605740 $Y=648220
X5047 584 1 2 591 3447 3470 1233 ICV_27 $T=619380 557880 1 0 $X=619380 $Y=552460
X5048 3360 1 3351 3384 2 ND2T $T=613800 628440 1 180 $X=608840 $Y=628060
X5049 3330 563 1 2 BUF6 $T=606360 578040 0 0 $X=606360 $Y=577660
X5050 237 221 2321 2299 2 1 MXL2HS $T=424700 547800 0 180 $X=419120 $Y=542380
X5051 238 221 2327 2307 2 1 MXL2HS $T=425320 557880 1 180 $X=419740 $Y=557500
X5052 2349 2260 2333 2014 2 1 MXL2HS $T=426560 578040 1 180 $X=420980 $Y=577660
X5053 3226 3216 3240 3254 2 1 MXL2HS $T=582180 658680 0 0 $X=582180 $Y=658300
X5054 2794 3212 3228 3245 1 2 HA1P $T=576600 688920 0 0 $X=576600 $Y=688540
X5055 1648 1 1672 1653 1690 1704 2 1648 1704 1653 113 1726 1233 ICV_28 $T=301940 557880 1 0 $X=301940 $Y=552460
X5056 1742 1 1763 1733 131 1790 2 1742 1790 1733 1800 1808 1233 ICV_28 $T=316200 547800 0 0 $X=316200 $Y=547420
X5057 1645 1 1761 1801 137 1795 2 1795 1727 1761 139 1807 1233 ICV_28 $T=321160 557880 0 0 $X=321160 $Y=557500
X5058 1919 1 1892 1908 170 1957 2 1973 1893 1978 175 1983 1233 ICV_28 $T=352160 547800 1 0 $X=352160 $Y=542380
X5059 1973 1 1983 1994 178 1978 2 1973 1994 1978 186 2030 1233 ICV_28 $T=360840 547800 1 0 $X=360840 $Y=542380
X5060 1975 1 1981 1876 181 2006 2 1975 2006 1876 2022 2023 1233 ICV_28 $T=361460 567960 1 0 $X=361460 $Y=562540
X5061 2127 1 2117 2041 2176 2120 2 2162 2120 2041 2189 2188 1233 ICV_28 $T=392460 557880 1 0 $X=392460 $Y=552460
X5062 2100 1 2109 2070 2192 2157 2 2100 2157 2204 2220 2070 1233 ICV_28 $T=395560 567960 0 0 $X=395560 $Y=567580
X5063 2642 1 2676 2696 2714 2713 2 2642 2696 2723 2740 2713 1233 ICV_28 $T=485460 658680 0 0 $X=485460 $Y=658300
X5064 2734 1 2746 2781 2751 2762 2 2734 2781 2774 2771 2762 1233 ICV_28 $T=496620 678840 0 0 $X=496620 $Y=678460
X5065 3094 1 3099 3101 3100 3107 2 3094 3101 3116 3119 3107 1233 ICV_28 $T=553660 618360 1 0 $X=553660 $Y=612940
X5066 1864 1925 1985 2 1 1940 XNR3 $T=350920 608280 0 0 $X=350920 $Y=607900
.ENDS
***************************************
.SUBCKT ANTENNA GND VCC A
** N=4 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 DELB $T=9920 0 0 0 $X=9920 $Y=-380
X1 5 2 3 6 7 8 9 ICV_4 $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT AN4B1 I3 I2 I1 O B1 GND VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF8CK I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN2S I1 I2 GND O VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV4 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MOAI1HP B2 B1 GND A1 O A2 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI22H B2 B1 GND A2 O A1 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNR2H I2 O I1 GND VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO112 O C2 C1 VCC B1 GND A1
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO222 C1 C2 B2 B1 A1 A2 GND VCC O
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA222S A2 A1 B2 B1 C2 C1 VCC GND O
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT QDFFRBS D CK RB VCC GND Q
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI12H B2 B1 VCC O A1 GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540
+ 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560
+ 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580
+ 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640
+ 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660
+ 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680
+ 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700
+ 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720
+ 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740
+ 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760
+ 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780
+ 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800
+ 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820
+ 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840
+ 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860
+ 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880
+ 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900
+ 901 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920
+ 921 922 923 924 925 926 927 928 929 930 931 932 933 934 935 936 937 938 939 940
+ 941 942 943 944 945 946 947 948 949 950 951 952 953 954 955 956 957 958 959 960
+ 961 962 963 964 965 966 967 968 969 970 971 972 973 974 975 976 977 978 979 980
+ 981 982 983 984 985 986 987 988 989 990 991 992 993 994 995 996 997 998 999 1000
+ 1001 1002 1003 1004 1005 1006 1007 1008 1009 1010 1011 1012 1013 1014 1015 1016 1017 1018 1019 1020
+ 1021 1022 1023 1024 1025 1026 1027 1028 1029 1030 1031 1032 1033 1034 1035 1036 1037 1038 1039 1040
+ 1041 1042 1043 1044 1045 1046 1047 1048 1049 1050 1051 1052 1053 1054 1055 1056 1057 1058 1059 1060
+ 1061 1062 1063 1064 1065 1066 1067 1068 1069 1070 1071 1072 1073 1074 1075 1076 1077 1078 1079 1080
+ 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 1093 1094 1095 1096 1097 1098 1099 1100
+ 1101 1102 1103 1104 1105 1106 1107 1108 1109 1110 1111 1112 1113 1114 1115 1116 1117 1118 1119 1120
+ 1121 1122 1123 1124 1125 1126 1127 1128 1129 1130 1131 1132 1133 1134 1135 1136 1137 1138 1139 1156
+ 1202
** N=6144 EP=1141 IP=31563 FDC=0
X0 1138 6141 6141 6141 1156 6141 1139 YA2GSD $T=1349740 417270 0 90 $X=1210240 $Y=420120
X1 1215 2 1203 1 INV1S $T=221960 436920 1 180 $X=220720 $Y=436540
X2 1204 2 1221 1 INV1S $T=220720 447000 0 0 $X=220720 $Y=446620
X3 1210 2 1220 1 INV1S $T=221960 527640 0 0 $X=221960 $Y=527260
X4 1216 2 1222 1 INV1S $T=222580 406680 0 0 $X=222580 $Y=406300
X5 1218 2 1226 1 INV1S $T=223200 376440 0 0 $X=223200 $Y=376060
X6 1225 2 1237 1 INV1S $T=225060 396600 1 0 $X=225060 $Y=391180
X7 1232 2 1240 1 INV1S $T=225680 467160 0 0 $X=225680 $Y=466780
X8 1209 2 1228 1 INV1S $T=228160 517560 1 180 $X=226920 $Y=517180
X9 1208 2 1262 1 INV1S $T=230020 447000 0 0 $X=230020 $Y=446620
X10 1206 2 1267 1 INV1S $T=230640 386520 1 0 $X=230640 $Y=381100
X11 1259 2 1231 1 INV1S $T=230640 467160 0 0 $X=230640 $Y=466780
X12 1262 2 1269 1 INV1S $T=231260 447000 1 0 $X=231260 $Y=441580
X13 1288 2 1296 1 INV1S $T=236220 497400 0 0 $X=236220 $Y=497020
X14 1250 2 1331 1 INV1S $T=240560 527640 1 0 $X=240560 $Y=522220
X15 1262 2 1348 1 INV1S $T=244280 447000 1 0 $X=244280 $Y=441580
X16 1264 2 1316 1 INV1S $T=245520 477240 1 180 $X=244280 $Y=476860
X17 49 2 35 1 INV1S $T=249860 497400 1 180 $X=248620 $Y=497020
X18 1267 2 1343 1 INV1S $T=251720 386520 1 0 $X=251720 $Y=381100
X19 1267 2 1413 1 INV1S $T=257300 386520 1 0 $X=257300 $Y=381100
X20 1403 2 1392 1 INV1S $T=257920 517560 1 0 $X=257920 $Y=512140
X21 1383 2 1395 1 INV1S $T=258540 527640 0 0 $X=258540 $Y=527260
X22 1353 2 1414 1 INV1S $T=260400 406680 1 0 $X=260400 $Y=401260
X23 1413 2 1433 1 INV1S $T=265980 386520 1 0 $X=265980 $Y=381100
X24 1420 2 1458 1 INV1S $T=270940 517560 0 0 $X=270940 $Y=517180
X25 70 2 1481 1 INV1S $T=274040 527640 0 0 $X=274040 $Y=527260
X26 1590 2 1612 1 INV1S $T=296980 386520 1 0 $X=296980 $Y=381100
X27 1602 2 1620 1 INV1S $T=298220 376440 1 0 $X=298220 $Y=371020
X28 1610 2 1626 1 INV1S $T=300080 396600 1 0 $X=300080 $Y=391180
X29 1591 2 1636 1 INV1S $T=301320 376440 0 0 $X=301320 $Y=376060
X30 1684 2 1534 1 INV1S $T=302560 467160 0 180 $X=301320 $Y=461740
X31 1635 2 1660 1 INV1S $T=303800 396600 1 0 $X=303800 $Y=391180
X32 1629 2 1675 1 INV1S $T=303800 447000 0 0 $X=303800 $Y=446620
X33 1667 2 1680 1 INV1S $T=306280 406680 1 0 $X=306280 $Y=401260
X34 1665 2 1677 1 INV1S $T=306280 436920 0 0 $X=306280 $Y=436540
X35 1649 2 1671 1 INV1S $T=308140 447000 1 180 $X=306900 $Y=446620
X36 1634 2 1703 1 INV1S $T=308760 366360 0 0 $X=308760 $Y=365980
X37 1689 2 1704 1 INV1S $T=308760 396600 0 0 $X=308760 $Y=396220
X38 1638 2 1705 1 INV1S $T=308760 426840 1 0 $X=308760 $Y=421420
X39 1651 2 1716 1 INV1S $T=309380 376440 0 0 $X=309380 $Y=376060
X40 1710 2 1702 1 INV1S $T=311240 396600 1 180 $X=310000 $Y=396220
X41 1712 2 1699 1 INV1S $T=310000 457080 1 0 $X=310000 $Y=451660
X42 1684 2 1727 1 INV1S $T=310000 467160 0 0 $X=310000 $Y=466780
X43 1694 2 1734 1 INV1S $T=310000 487320 1 0 $X=310000 $Y=481900
X44 1674 2 1684 1 INV1S $T=311240 497400 1 180 $X=310000 $Y=497020
X45 92 2 1719 1 INV1S $T=310620 366360 0 0 $X=310620 $Y=365980
X46 1751 2 1718 1 INV1S $T=312480 497400 0 180 $X=311240 $Y=491980
X47 1607 2 1737 1 INV1S $T=312480 386520 0 0 $X=312480 $Y=386140
X48 1623 2 1761 1 INV1S $T=313720 436920 1 0 $X=313720 $Y=431500
X49 1759 2 1731 1 INV1S $T=316200 497400 0 0 $X=316200 $Y=497020
X50 1778 2 1746 1 INV1S $T=319920 497400 1 180 $X=318680 $Y=497020
X51 109 2 1789 1 INV1S $T=319300 537720 1 0 $X=319300 $Y=532300
X52 1687 2 1768 1 INV1S $T=320540 497400 1 0 $X=320540 $Y=491980
X53 1797 2 1784 1 INV1S $T=321780 497400 1 180 $X=320540 $Y=497020
X54 129 2 1871 1 INV1S $T=340380 386520 0 180 $X=339140 $Y=381100
X55 1891 2 1917 1 INV1S $T=341620 507480 0 0 $X=341620 $Y=507100
X56 1815 2 1911 1 INV1S $T=344720 386520 0 0 $X=344720 $Y=386140
X57 1845 2 1933 1 INV1S $T=347820 386520 0 0 $X=347820 $Y=386140
X58 1914 2 1979 1 INV1S $T=354640 366360 0 0 $X=354640 $Y=365980
X59 1960 2 1990 1 INV1S $T=355880 386520 1 0 $X=355880 $Y=381100
X60 2014 2 2019 1 INV1S $T=362700 507480 0 0 $X=362700 $Y=507100
X61 2029 2 1949 1 INV1S $T=363940 517560 0 180 $X=362700 $Y=512140
X62 2070 2 2003 1 INV1S $T=369520 507480 1 180 $X=368280 $Y=507100
X63 162 2 2062 1 INV1S $T=368900 477240 0 0 $X=368900 $Y=476860
X64 2070 2 1835 1 INV1S $T=368900 507480 1 0 $X=368900 $Y=502060
X65 2080 2 2070 1 INV1S $T=370760 507480 1 180 $X=369520 $Y=507100
X66 1840 2 2095 1 INV1S $T=370760 376440 0 0 $X=370760 $Y=376060
X67 167 2 2130 1 INV1S $T=378820 487320 0 180 $X=377580 $Y=481900
X68 2168 2 2096 1 INV1S $T=383780 447000 1 180 $X=382540 $Y=446620
X69 154 2 2182 1 INV1S $T=384400 487320 0 0 $X=384400 $Y=486940
X70 2202 2 2213 1 INV1S $T=389360 507480 0 0 $X=389360 $Y=507100
X71 180 2 2091 1 INV1S $T=392460 447000 0 180 $X=391220 $Y=441580
X72 181 2 2194 1 INV1S $T=392460 487320 1 180 $X=391220 $Y=486940
X73 173 2 2216 1 INV1S $T=392460 457080 1 0 $X=392460 $Y=451660
X74 2130 2 2227 1 INV1S $T=392460 457080 0 0 $X=392460 $Y=456700
X75 2227 2 2186 1 INV1S $T=394320 447000 0 180 $X=393080 $Y=441580
X76 194 2 2046 1 INV1S $T=396180 447000 0 180 $X=394940 $Y=441580
X77 2227 2 2236 1 INV1S $T=394940 447000 0 0 $X=394940 $Y=446620
X78 166 2 2225 1 INV1S $T=398660 416760 0 180 $X=397420 $Y=411340
X79 2245 2 2168 1 INV1S $T=398660 457080 0 180 $X=397420 $Y=451660
X80 192 2 2184 1 INV1S $T=398660 497400 1 180 $X=397420 $Y=497020
X81 2246 2 2271 1 INV1S $T=399280 507480 1 0 $X=399280 $Y=502060
X82 197 2 2268 1 INV1S $T=401140 467160 1 180 $X=399900 $Y=466780
X83 2268 2 2198 1 INV1S $T=401760 436920 1 180 $X=400520 $Y=436540
X84 193 2 2280 1 INV1S $T=400520 497400 1 0 $X=400520 $Y=491980
X85 2270 2 2256 1 INV1S $T=401760 507480 1 180 $X=400520 $Y=507100
X86 2268 2 2061 1 INV1S $T=401140 457080 0 0 $X=401140 $Y=456700
X87 199 2 195 1 INV1S $T=402380 376440 0 0 $X=402380 $Y=376060
X88 202 2 2260 1 INV1S $T=403620 447000 0 180 $X=402380 $Y=441580
X89 201 2 2288 1 INV1S $T=403000 386520 1 0 $X=403000 $Y=381100
X90 201 2 2149 1 INV1S $T=403000 426840 1 0 $X=403000 $Y=421420
X91 162 2 2317 1 INV1S $T=406100 477240 1 0 $X=406100 $Y=471820
X92 2344 2 2282 1 INV1S $T=412300 477240 1 180 $X=411060 $Y=476860
X93 193 2 2347 1 INV1S $T=411060 507480 1 0 $X=411060 $Y=502060
X94 210 2 2344 1 INV1S $T=414780 487320 0 180 $X=413540 $Y=481900
X95 2412 2 2416 1 INV1S $T=425320 497400 0 0 $X=425320 $Y=497020
X96 2415 2 2414 1 INV1S $T=427800 426840 1 180 $X=426560 $Y=426460
X97 2417 2 2430 1 INV1S $T=427800 507480 1 0 $X=427800 $Y=502060
X98 229 2 2420 1 INV1S $T=428420 376440 0 0 $X=428420 $Y=376060
X99 232 2 2421 1 INV1S $T=433380 426840 0 180 $X=432140 $Y=421420
X100 135 2 2465 1 INV1S $T=434000 447000 1 0 $X=434000 $Y=441580
X101 2212 2 2467 1 INV1S $T=434620 447000 0 0 $X=434620 $Y=446620
X102 2468 2 2446 1 INV1S $T=435860 507480 0 180 $X=434620 $Y=502060
X103 2467 2 215 1 INV1S $T=437720 366360 1 180 $X=436480 $Y=365980
X104 243 2 238 1 INV1S $T=438960 537720 0 180 $X=437720 $Y=532300
X105 2454 2 2492 1 INV1S $T=438340 517560 1 0 $X=438340 $Y=512140
X106 2450 2 2511 1 INV1S $T=438960 527640 1 0 $X=438960 $Y=522220
X107 2501 2 2433 1 INV1S $T=440820 477240 0 180 $X=439580 $Y=471820
X108 2500 2 2505 1 INV1S $T=440200 457080 1 0 $X=440200 $Y=451660
X109 234 2 2530 1 INV1S $T=441440 426840 0 0 $X=441440 $Y=426460
X110 2469 2 2514 1 INV1S $T=443300 527640 0 180 $X=442060 $Y=522220
X111 2536 2 2523 1 INV1S $T=445780 487320 1 180 $X=444540 $Y=486940
X112 256 2 2501 1 INV1S $T=447640 497400 1 180 $X=446400 $Y=497020
X113 2501 2 2488 1 INV1S $T=447020 487320 1 0 $X=447020 $Y=481900
X114 2554 2 2529 1 INV1S $T=448880 436920 1 180 $X=447640 $Y=436540
X115 2520 2 2537 1 INV1S $T=447640 447000 0 0 $X=447640 $Y=446620
X116 2557 2 2544 1 INV1S $T=449500 467160 1 180 $X=448260 $Y=466780
X117 235 2 2556 1 INV1S $T=450120 436920 1 0 $X=450120 $Y=431500
X118 2573 2 2558 1 INV1S $T=451980 426840 0 180 $X=450740 $Y=421420
X119 260 2 262 1 INV1S $T=453220 376440 1 0 $X=453220 $Y=371020
X120 2589 2 2590 1 INV1S $T=455080 426840 0 0 $X=455080 $Y=426460
X121 2584 2 193 1 INV1S $T=455080 497400 1 0 $X=455080 $Y=491980
X122 2613 2 2604 1 INV1S $T=459420 497400 1 0 $X=459420 $Y=491980
X123 2380 2 270 1 INV1S $T=463140 376440 0 0 $X=463140 $Y=376060
X124 2576 2 2632 1 INV1S $T=464380 396600 0 180 $X=463140 $Y=391180
X125 2617 2 2630 1 INV1S $T=465000 487320 0 180 $X=463760 $Y=481900
X126 272 2 2656 1 INV1S $T=465620 376440 0 0 $X=465620 $Y=376060
X127 275 2 264 1 INV1S $T=467480 366360 1 180 $X=466240 $Y=365980
X128 2372 2 275 1 INV1S $T=466240 416760 0 0 $X=466240 $Y=416380
X129 2516 2 2695 1 INV1S $T=468720 497400 1 0 $X=468720 $Y=491980
X130 2685 2 273 1 INV1S $T=471200 416760 1 180 $X=469960 $Y=416380
X131 2574 2 2687 1 INV1S $T=469960 426840 1 0 $X=469960 $Y=421420
X132 2399 2 240 1 INV1S $T=470580 396600 1 0 $X=470580 $Y=391180
X133 2611 2 2698 1 INV1S $T=470580 487320 0 0 $X=470580 $Y=486940
X134 246 2 290 1 INV1S $T=471820 386520 1 0 $X=471820 $Y=381100
X135 2727 2 272 1 INV1S $T=474920 426840 1 180 $X=473680 $Y=426460
X136 2605 2 2707 1 INV1S $T=473680 497400 1 0 $X=473680 $Y=491980
X137 2485 2 2680 1 INV1S $T=475540 406680 0 0 $X=475540 $Y=406300
X138 2684 2 2731 1 INV1S $T=479880 477240 1 180 $X=478640 $Y=476860
X139 2675 2 2737 1 INV1S $T=478640 487320 0 0 $X=478640 $Y=486940
X140 2739 2 2631 1 INV1S $T=479880 497400 0 180 $X=478640 $Y=491980
X141 2606 2 2746 1 INV1S $T=478640 497400 0 0 $X=478640 $Y=497020
X142 2748 2 2739 1 INV1S $T=481120 477240 1 180 $X=479880 $Y=476860
X143 2739 2 295 1 INV1S $T=480500 497400 1 0 $X=480500 $Y=491980
X144 296 2 276 1 INV1S $T=482360 537720 0 180 $X=481120 $Y=532300
X145 225 2 2533 1 INV1S $T=481740 396600 1 0 $X=481740 $Y=391180
X146 2585 2 2555 1 INV1S $T=483600 457080 1 180 $X=482360 $Y=456700
X147 2760 2 296 1 INV1S $T=483600 497400 0 180 $X=482360 $Y=491980
X148 303 2 278 1 INV1S $T=483600 517560 0 180 $X=482360 $Y=512140
X149 2773 2 301 1 INV1S $T=485460 386520 0 180 $X=484220 $Y=381100
X150 312 2 308 1 INV1S $T=487940 537720 0 180 $X=486700 $Y=532300
X151 2786 2 2797 1 INV1S $T=487940 376440 0 0 $X=487940 $Y=376060
X152 2763 2 2621 1 INV1S $T=487940 416760 1 0 $X=487940 $Y=411340
X153 315 2 2659 1 INV1S $T=489180 517560 1 180 $X=487940 $Y=517180
X154 2795 2 315 1 INV1S $T=490420 507480 1 180 $X=489180 $Y=507100
X155 2814 2 303 1 INV1S $T=492900 497400 1 180 $X=491660 $Y=497020
X156 131 2 323 1 INV1S $T=493520 376440 1 0 $X=493520 $Y=371020
X157 2826 2 2795 1 INV1S $T=494760 497400 1 180 $X=493520 $Y=497020
X158 2815 2 2842 1 INV1S $T=494760 406680 1 0 $X=494760 $Y=401260
X159 2838 2 2760 1 INV1S $T=496620 487320 1 180 $X=495380 $Y=486940
X160 2800 2 2802 1 INV1S $T=496000 396600 0 0 $X=496000 $Y=396220
X161 2809 2 2730 1 INV1S $T=496620 436920 1 0 $X=496620 $Y=431500
X162 2851 2 2814 1 INV1S $T=497860 497400 0 180 $X=496620 $Y=491980
X163 2856 2 2862 1 INV1S $T=497860 447000 0 0 $X=497860 $Y=446620
X164 2854 2 2863 1 INV1S $T=498480 447000 1 0 $X=498480 $Y=441580
X165 2870 2 2705 1 INV1S $T=500340 416760 0 180 $X=499100 $Y=411340
X166 2860 2 2866 1 INV1S $T=502200 447000 0 180 $X=500960 $Y=441580
X167 2858 2 2890 1 INV1S $T=501580 507480 1 0 $X=501580 $Y=502060
X168 2888 2 2861 1 INV1S $T=503440 406680 1 180 $X=502200 $Y=406300
X169 2811 2 2880 1 INV1S $T=502200 416760 0 0 $X=502200 $Y=416380
X170 2796 2 2899 1 INV1S $T=502200 507480 0 0 $X=502200 $Y=507100
X171 324 2 2891 1 INV1S $T=502200 517560 0 0 $X=502200 $Y=517180
X172 2885 2 328 1 INV1S $T=504060 527640 0 0 $X=504060 $Y=527260
X173 2842 2 2836 1 INV1S $T=505920 406680 0 180 $X=504680 $Y=401260
X174 2901 2 2875 1 INV1S $T=505920 416760 1 180 $X=504680 $Y=416380
X175 2908 2 2887 1 INV1S $T=505920 436920 1 180 $X=504680 $Y=436540
X176 2909 2 317 1 INV1S $T=506540 527640 1 180 $X=505300 $Y=527260
X177 2888 2 2905 1 INV1S $T=506540 406680 0 0 $X=506540 $Y=406300
X178 2906 2 2888 1 INV1S $T=507780 416760 1 180 $X=506540 $Y=416380
X179 2834 2 2753 1 INV1S $T=506540 426840 1 0 $X=506540 $Y=421420
X180 2900 2 2915 1 INV1S $T=506540 436920 0 0 $X=506540 $Y=436540
X181 2911 2 300 1 INV1S $T=507780 527640 1 180 $X=506540 $Y=527260
X182 2928 2 333 1 INV1S $T=509020 527640 1 180 $X=507780 $Y=527260
X183 2935 2 2920 1 INV1S $T=509640 416760 0 180 $X=508400 $Y=411340
X184 2934 2 336 1 INV1S $T=509020 537720 1 0 $X=509020 $Y=532300
X185 2922 2 2897 1 INV1S $T=509640 447000 1 0 $X=509640 $Y=441580
X186 2945 2 2955 1 INV1S $T=511500 436920 1 0 $X=511500 $Y=431500
X187 2467 2 2966 1 INV1S $T=512740 436920 0 0 $X=512740 $Y=436540
X188 2949 2 2961 1 INV1S $T=512740 447000 1 0 $X=512740 $Y=441580
X189 2967 2 2964 1 INV1S $T=513980 447000 1 180 $X=512740 $Y=446620
X190 2855 2 2729 1 INV1S $T=513360 436920 1 0 $X=513360 $Y=431500
X191 2667 2 2989 1 INV1S $T=514600 447000 0 0 $X=514600 $Y=446620
X192 2916 2 304 1 INV1S $T=514600 527640 1 0 $X=514600 $Y=522220
X193 2988 2 3001 1 INV1S $T=515840 406680 0 0 $X=515840 $Y=406300
X194 2998 2 3003 1 INV1S $T=515840 426840 0 0 $X=515840 $Y=426460
X195 2989 2 3006 1 INV1S $T=515840 447000 1 0 $X=515840 $Y=441580
X196 3010 2 2981 1 INV1S $T=517700 457080 0 180 $X=516460 $Y=451660
X197 3007 2 3015 1 INV1S $T=517080 386520 0 0 $X=517080 $Y=386140
X198 3051 2 3016 1 INV1S $T=518940 447000 1 180 $X=517700 $Y=446620
X199 3007 2 344 1 INV1S $T=518320 376440 1 0 $X=518320 $Y=371020
X200 2993 2 3007 1 INV1S $T=519560 406680 1 180 $X=518320 $Y=406300
X201 3031 2 3027 1 INV1S $T=520800 457080 0 180 $X=519560 $Y=451660
X202 3046 2 302 1 INV1S $T=523280 537720 0 180 $X=522040 $Y=532300
X203 3035 2 3063 1 INV1S $T=523280 416760 0 0 $X=523280 $Y=416380
X204 2939 2 3088 1 INV1S $T=523280 447000 1 0 $X=523280 $Y=441580
X205 3061 2 3075 1 INV1S $T=523900 436920 1 0 $X=523900 $Y=431500
X206 2771 2 3092 1 INV1S $T=525140 487320 1 0 $X=525140 $Y=481900
X207 3074 2 3009 1 INV1S $T=527000 436920 0 180 $X=525760 $Y=431500
X208 2879 2 3123 1 INV1S $T=529480 376440 0 0 $X=529480 $Y=376060
X209 3093 2 3122 1 INV1S $T=530100 507480 0 0 $X=530100 $Y=507100
X210 3139 2 3066 1 INV1S $T=531960 376440 1 180 $X=530720 $Y=376060
X211 3002 2 3139 1 INV1S $T=530720 396600 0 0 $X=530720 $Y=396220
X212 3128 2 3130 1 INV1S $T=530720 436920 1 0 $X=530720 $Y=431500
X213 2812 2 3137 1 INV1S $T=530720 497400 0 0 $X=530720 $Y=497020
X214 3081 2 3162 1 INV1S $T=532580 487320 0 0 $X=532580 $Y=486940
X215 3153 2 3047 1 INV1S $T=534440 436920 0 180 $X=533200 $Y=431500
X216 3163 2 3038 1 INV1S $T=535680 436920 0 180 $X=534440 $Y=431500
X217 3157 2 3168 1 INV1S $T=535680 396600 1 0 $X=535680 $Y=391180
X218 3162 2 3113 1 INV1S $T=537540 477240 1 180 $X=536300 $Y=476860
X219 3162 2 3175 1 INV1S $T=536300 497400 1 0 $X=536300 $Y=491980
X220 2932 2 3131 1 INV1S $T=537540 447000 1 0 $X=537540 $Y=441580
X221 3190 2 3106 1 INV1S $T=539400 416760 0 180 $X=538160 $Y=411340
X222 3139 2 383 1 INV1S $T=538780 386520 1 0 $X=538780 $Y=381100
X223 385 2 3198 1 INV1S $T=541880 396600 1 180 $X=540640 $Y=396220
X224 3180 2 3233 1 INV1S $T=546220 416760 0 0 $X=546220 $Y=416380
X225 3238 2 3257 1 INV1S $T=548700 396600 1 0 $X=548700 $Y=391180
X226 341 2 2837 1 INV1S $T=551180 426840 1 180 $X=549940 $Y=426460
X227 3119 2 3266 1 INV1S $T=551800 487320 1 180 $X=550560 $Y=486940
X228 2948 2 3269 1 INV1S $T=553040 406680 0 180 $X=551800 $Y=401260
X229 400 2 3240 1 INV1S $T=553040 527640 1 180 $X=551800 $Y=527260
X230 366 2 3275 1 INV1S $T=553660 376440 0 180 $X=552420 $Y=371020
X231 3273 2 3278 1 INV1S $T=553660 416760 1 180 $X=552420 $Y=416380
X232 3175 2 3285 1 INV1S $T=553040 487320 0 0 $X=553040 $Y=486940
X233 3297 2 3292 1 INV1S $T=555520 416760 1 180 $X=554280 $Y=416380
X234 400 2 3288 1 INV1S $T=554900 527640 0 0 $X=554900 $Y=527260
X235 3223 2 3309 1 INV1S $T=555520 477240 0 0 $X=555520 $Y=476860
X236 2830 2 3314 1 INV1S $T=558000 467160 0 0 $X=558000 $Y=466780
X237 2992 2 3320 1 INV1S $T=559860 386520 1 180 $X=558620 $Y=386140
X238 3133 2 3313 1 INV1S $T=561100 386520 1 180 $X=559860 $Y=386140
X239 3331 2 3322 1 INV1S $T=561100 416760 1 180 $X=559860 $Y=416380
X240 3324 2 3316 1 INV1S $T=563580 406680 1 180 $X=562340 $Y=406300
X241 3349 2 3025 1 INV1S $T=565440 497400 1 180 $X=564200 $Y=497020
X242 3368 2 3373 1 INV1S $T=567300 497400 0 0 $X=567300 $Y=497020
X243 416 2 2941 1 INV1S $T=569160 507480 0 0 $X=569160 $Y=507100
X244 3287 2 423 1 INV1S $T=572880 487320 1 0 $X=572880 $Y=481900
X245 3253 2 3413 1 INV1S $T=574740 406680 0 0 $X=574740 $Y=406300
X246 423 2 3020 1 INV1S $T=576600 487320 1 180 $X=575360 $Y=486940
X247 3297 2 3276 1 INV1S $T=577220 386520 0 180 $X=575980 $Y=381100
X248 3426 2 3424 1 INV1S $T=577840 376440 0 180 $X=576600 $Y=371020
X249 431 2 435 1 INV1S $T=579700 366360 0 0 $X=579700 $Y=365980
X250 441 2 3476 1 INV1S $T=587140 376440 0 180 $X=585900 $Y=371020
X251 3445 2 3471 1 INV1S $T=587760 386520 1 180 $X=586520 $Y=386140
X252 3442 2 3507 1 INV1S $T=587140 376440 0 0 $X=587140 $Y=376060
X253 3495 2 3511 1 INV1S $T=589620 396600 1 0 $X=589620 $Y=391180
X254 3505 2 3510 1 INV1S $T=589620 416760 0 0 $X=589620 $Y=416380
X255 3520 2 3530 1 INV1S $T=592100 386520 0 0 $X=592100 $Y=386140
X256 3524 2 3529 1 INV1S $T=592720 416760 0 0 $X=592720 $Y=416380
X257 3431 2 3492 1 INV1S $T=595820 386520 0 180 $X=594580 $Y=381100
X258 3536 2 3527 1 INV1S $T=595820 396600 0 180 $X=594580 $Y=391180
X259 3526 2 3532 1 INV1S $T=597060 436920 1 0 $X=597060 $Y=431500
X260 3549 2 3525 1 INV1S $T=598920 416760 0 180 $X=597680 $Y=411340
X261 3566 2 3540 1 INV1S $T=600160 416760 0 180 $X=598920 $Y=411340
X262 3581 2 3428 1 INV1S $T=600780 436920 0 180 $X=599540 $Y=431500
X263 3563 2 3573 1 INV1S $T=600160 416760 0 0 $X=600160 $Y=416380
X264 3568 2 3547 1 INV1S $T=600160 426840 1 0 $X=600160 $Y=421420
X265 405 2 3557 1 INV1S $T=602640 477240 0 180 $X=601400 $Y=471820
X266 439 2 3591 1 INV1S $T=603260 366360 0 0 $X=603260 $Y=365980
X267 3613 2 3595 1 INV1S $T=608840 416760 1 180 $X=607600 $Y=416380
X268 3537 2 3619 1 INV1S $T=607600 426840 1 0 $X=607600 $Y=421420
X269 3606 2 3631 1 INV1S $T=613180 436920 0 180 $X=611940 $Y=431500
X270 3657 2 3569 1 INV1S $T=614420 436920 0 180 $X=613180 $Y=431500
X271 3671 2 3665 1 INV1S $T=615660 426840 1 180 $X=614420 $Y=426460
X272 3545 2 3694 1 INV1S $T=617520 507480 0 0 $X=617520 $Y=507100
X273 3730 2 3680 1 INV1S $T=624340 396600 1 180 $X=623100 $Y=396220
X274 3493 2 3738 1 INV1S $T=624340 406680 1 0 $X=624340 $Y=401260
X275 3730 2 3754 1 INV1S $T=628060 406680 1 0 $X=628060 $Y=401260
X276 3601 2 3778 1 INV1S $T=629920 497400 0 0 $X=629920 $Y=497020
X277 3601 2 3771 1 INV1S $T=631160 507480 1 0 $X=631160 $Y=502060
X278 473 2 3796 1 INV1S $T=634880 376440 1 0 $X=634880 $Y=371020
X279 3833 2 3831 1 INV1S $T=644800 406680 1 180 $X=643560 $Y=406300
X280 3421 2 3855 1 INV1S $T=644800 416760 0 0 $X=644800 $Y=416380
X281 3443 2 3891 1 INV1S $T=652240 386520 0 0 $X=652240 $Y=386140
X282 3895 2 3881 1 INV1S $T=654100 396600 1 180 $X=652860 $Y=396220
X283 513 2 3930 1 INV1S $T=657200 527640 1 0 $X=657200 $Y=522220
X284 3930 2 3948 1 INV1S $T=659680 507480 1 0 $X=659680 $Y=502060
X285 3942 2 3921 1 INV1S $T=660300 447000 0 0 $X=660300 $Y=446620
X286 510 2 3953 1 INV1S $T=662780 366360 1 180 $X=661540 $Y=365980
X287 3953 2 511 1 INV1S $T=662160 376440 1 0 $X=662160 $Y=371020
X288 3930 2 3972 1 INV1S $T=663400 527640 0 0 $X=663400 $Y=527260
X289 4071 2 3971 1 INV1S $T=684480 497400 0 180 $X=683240 $Y=491980
X290 4071 2 4073 1 INV1S $T=684480 497400 1 0 $X=684480 $Y=491980
X291 545 2 4071 1 INV1S $T=686340 507480 1 180 $X=685100 $Y=507100
X292 2465 2 4136 1 INV1S $T=705560 426840 1 180 $X=704320 $Y=426460
X293 4219 2 4192 1 INV1S $T=716100 396600 0 180 $X=714860 $Y=391180
X294 4336 2 4239 1 INV1S $T=738420 416760 0 0 $X=738420 $Y=416380
X295 604 2 564 1 INV1S $T=738420 537720 1 0 $X=738420 $Y=532300
X296 606 2 4210 1 INV1S $T=740900 447000 0 180 $X=739660 $Y=441580
X297 4354 2 4324 1 INV1S $T=743380 457080 1 0 $X=743380 $Y=451660
X298 4368 2 4348 1 INV1S $T=746480 467160 1 180 $X=745240 $Y=466780
X299 4372 2 4188 1 INV1S $T=746480 477240 0 180 $X=745240 $Y=471820
X300 4363 2 4276 1 INV1S $T=745240 517560 0 0 $X=745240 $Y=517180
X301 4365 2 4220 1 INV1S $T=745860 457080 1 0 $X=745860 $Y=451660
X302 4188 2 4368 1 INV1S $T=746480 467160 0 0 $X=746480 $Y=466780
X303 4371 2 3995 1 INV1S $T=747100 497400 1 0 $X=747100 $Y=491980
X304 4380 2 4205 1 INV1S $T=748960 467160 1 180 $X=747720 $Y=466780
X305 4389 2 4197 1 INV1S $T=750200 497400 0 180 $X=748960 $Y=491980
X306 4387 2 4173 1 INV1S $T=750200 527640 1 180 $X=748960 $Y=527260
X307 622 2 4390 1 INV1S $T=750820 517560 1 180 $X=749580 $Y=517180
X308 4392 2 4322 1 INV1S $T=751440 386520 0 180 $X=750200 $Y=381100
X309 4398 2 4152 1 INV1S $T=752060 396600 0 0 $X=752060 $Y=396220
X310 4402 2 4268 1 INV1S $T=755160 426840 1 0 $X=755160 $Y=421420
X311 4368 2 4416 1 INV1S $T=755160 467160 0 0 $X=755160 $Y=466780
X312 4418 2 4377 1 INV1S $T=757020 436920 0 180 $X=755780 $Y=431500
X313 4418 2 4303 1 INV1S $T=757020 436920 1 180 $X=755780 $Y=436540
X314 632 2 626 1 INV1S $T=757020 537720 0 180 $X=755780 $Y=532300
X315 4404 2 4418 1 INV1S $T=757640 447000 0 180 $X=756400 $Y=441580
X316 4338 2 4438 1 INV1S $T=759500 497400 0 0 $X=759500 $Y=497020
X317 4438 2 4252 1 INV1S $T=763220 497400 1 180 $X=761980 $Y=497020
X318 632 2 4216 1 INV1S $T=764460 497400 1 180 $X=763220 $Y=497020
X319 632 2 4475 1 INV1S $T=765080 517560 0 0 $X=765080 $Y=517180
X320 632 2 4433 1 INV1S $T=766320 457080 1 0 $X=766320 $Y=451660
X321 4446 2 4408 1 INV1S $T=766940 396600 1 0 $X=766940 $Y=391180
X322 4438 2 4494 1 INV1S $T=770660 497400 0 0 $X=770660 $Y=497020
X323 4438 2 4483 1 INV1S $T=770660 507480 1 0 $X=770660 $Y=502060
X324 4508 2 4507 1 INV1S $T=773140 436920 0 0 $X=773140 $Y=436540
X325 645 2 4508 1 INV1S $T=773140 477240 1 0 $X=773140 $Y=471820
X326 4508 2 649 1 INV1S $T=775620 447000 1 0 $X=775620 $Y=441580
X327 4555 2 656 1 INV1S $T=784920 406680 1 180 $X=783680 $Y=406300
X328 4555 2 4597 1 INV1S $T=794840 406680 0 0 $X=794840 $Y=406300
X329 4555 2 4617 1 INV1S $T=798560 467160 0 0 $X=798560 $Y=466780
X330 4518 2 4628 1 INV1S $T=801040 376440 0 0 $X=801040 $Y=376060
X331 4555 2 4611 1 INV1S $T=801660 477240 1 0 $X=801660 $Y=471820
X332 4641 2 4436 1 INV1S $T=804140 487320 1 180 $X=802900 $Y=486940
X333 4628 2 684 1 INV1S $T=807860 376440 0 0 $X=807860 $Y=376060
X334 4555 2 4666 1 INV1S $T=808480 487320 0 0 $X=808480 $Y=486940
X335 4641 2 4682 1 INV1S $T=810960 487320 1 0 $X=810960 $Y=481900
X336 680 2 4641 1 INV1S $T=812820 527640 1 0 $X=812820 $Y=522220
X337 4712 2 4570 1 INV1S $T=817160 426840 0 180 $X=815920 $Y=421420
X338 591 2 4712 1 INV1S $T=817780 416760 0 0 $X=817780 $Y=416380
X339 4712 2 4717 1 INV1S $T=819640 426840 1 0 $X=819640 $Y=421420
X340 2465 2 4704 1 INV1S $T=826460 447000 1 0 $X=826460 $Y=441580
X341 4746 2 4752 1 INV1S $T=829560 467160 0 0 $X=829560 $Y=466780
X342 4762 2 4754 1 INV1S $T=833280 426840 0 0 $X=833280 $Y=426460
X343 4774 2 4779 1 INV1S $T=835140 426840 0 0 $X=835140 $Y=426460
X344 4755 2 4781 1 INV1S $T=836380 507480 1 0 $X=836380 $Y=502060
X345 4799 2 4793 1 INV1S $T=838860 396600 1 180 $X=837620 $Y=396220
X346 4797 2 4799 1 INV1S $T=840100 406680 0 180 $X=838860 $Y=401260
X347 4907 2 4849 1 INV1S $T=861800 376440 0 180 $X=860560 $Y=371020
X348 4910 2 4903 1 INV1S $T=861800 467160 1 180 $X=860560 $Y=466780
X349 736 2 4910 1 INV1S $T=860560 487320 1 0 $X=860560 $Y=481900
X350 4822 2 4932 1 INV1S $T=860560 507480 0 0 $X=860560 $Y=507100
X351 4918 2 4828 1 INV1S $T=862420 376440 1 180 $X=861180 $Y=376060
X352 4886 2 4907 1 INV1S $T=861800 396600 1 0 $X=861800 $Y=391180
X353 4916 2 4923 1 INV1S $T=863040 436920 0 0 $X=863040 $Y=436540
X354 4923 2 4918 1 INV1S $T=864280 416760 0 0 $X=864280 $Y=416380
X355 4907 2 4951 1 INV1S $T=866140 376440 1 0 $X=866140 $Y=371020
X356 4947 2 4928 1 INV1S $T=868000 426840 0 0 $X=868000 $Y=426460
X357 4918 2 783 1 INV1S $T=872960 376440 0 0 $X=872960 $Y=376060
X358 786 2 4988 1 INV1S $T=874820 537720 1 0 $X=874820 $Y=532300
X359 4988 2 4956 1 INV1S $T=877920 537720 0 180 $X=876680 $Y=532300
X360 4988 2 796 1 INV1S $T=878540 537720 1 0 $X=878540 $Y=532300
X361 5007 2 4971 1 INV1S $T=880400 477240 1 180 $X=879160 $Y=476860
X362 5019 2 791 1 INV1S $T=882880 396600 0 180 $X=881640 $Y=391180
X363 4955 2 5019 1 INV1S $T=882260 406680 1 0 $X=882260 $Y=401260
X364 4917 2 5050 1 INV1S $T=887840 467160 1 0 $X=887840 $Y=461740
X365 5054 2 5033 1 INV1S $T=890320 426840 1 180 $X=889080 $Y=426460
X366 5057 2 4964 1 INV1S $T=891560 477240 1 0 $X=891560 $Y=471820
X367 4781 2 5073 1 INV1S $T=892180 487320 1 0 $X=892180 $Y=481900
X368 5069 2 5014 1 INV1S $T=892800 426840 1 0 $X=892800 $Y=421420
X369 5073 2 5092 1 INV1S $T=894040 477240 0 0 $X=894040 $Y=476860
X370 5073 2 5082 1 INV1S $T=894660 487320 1 0 $X=894660 $Y=481900
X371 4932 2 5083 1 INV1S $T=896520 517560 0 180 $X=895280 $Y=512140
X372 5107 2 5038 1 INV1S $T=900860 517560 1 180 $X=899620 $Y=517180
X373 806 2 5107 1 INV1S $T=900860 527640 1 0 $X=900860 $Y=522220
X374 4932 2 5126 1 INV1S $T=903340 517560 1 0 $X=903340 $Y=512140
X375 5008 2 5155 1 INV1S $T=907680 467160 1 0 $X=907680 $Y=461740
X376 5155 2 5143 1 INV1S $T=908920 457080 1 0 $X=908920 $Y=451660
X377 5169 2 809 1 INV1S $T=910780 376440 1 180 $X=909540 $Y=376060
X378 5155 2 5163 1 INV1S $T=909540 467160 1 0 $X=909540 $Y=461740
X379 5081 2 5169 1 INV1S $T=912640 376440 1 180 $X=911400 $Y=376060
X380 5107 2 5179 1 INV1S $T=912640 517560 0 0 $X=912640 $Y=517180
X381 5169 2 836 1 INV1S $T=915740 376440 0 0 $X=915740 $Y=376060
X382 5201 2 5096 1 INV1S $T=918220 477240 0 0 $X=918220 $Y=476860
X383 5050 2 833 1 INV1S $T=925040 406680 1 180 $X=923800 $Y=406300
X384 5050 2 5240 1 INV1S $T=925040 406680 0 0 $X=925040 $Y=406300
X385 5278 2 5263 1 INV1S $T=933720 527640 0 180 $X=932480 $Y=522220
X386 860 2 830 1 INV1S $T=933100 497400 1 0 $X=933100 $Y=491980
X387 874 2 5278 1 INV1S $T=938060 537720 0 180 $X=936820 $Y=532300
X388 5323 2 5261 1 INV1S $T=944260 457080 0 180 $X=943020 $Y=451660
X389 5184 2 5323 1 INV1S $T=944260 457080 1 0 $X=944260 $Y=451660
X390 885 2 5184 1 INV1S $T=947360 436920 0 180 $X=946120 $Y=431500
X391 5323 2 5348 1 INV1S $T=948600 447000 0 0 $X=948600 $Y=446620
X392 5385 2 909 1 INV1S $T=958520 386520 0 0 $X=958520 $Y=386140
X393 860 2 5393 1 INV1S $T=961000 497400 1 0 $X=961000 $Y=491980
X394 5393 2 5412 1 INV1S $T=962240 497400 0 0 $X=962240 $Y=497020
X395 5412 2 924 1 INV1S $T=964100 517560 0 0 $X=964100 $Y=517180
X396 885 2 5364 1 INV1S $T=965340 426840 0 0 $X=965340 $Y=426460
X397 5440 2 5378 1 INV1S $T=974020 457080 0 0 $X=974020 $Y=456700
X398 5460 2 5427 1 INV1S $T=975880 477240 1 180 $X=974640 $Y=476860
X399 5412 2 931 1 INV1S $T=974640 507480 0 0 $X=974640 $Y=507100
X400 5455 2 942 1 INV1S $T=977740 376440 0 0 $X=977740 $Y=376060
X401 5376 2 5460 1 INV1S $T=977740 487320 1 0 $X=977740 $Y=481900
X402 924 2 5385 1 INV1S $T=980220 386520 0 0 $X=980220 $Y=386140
X403 5385 2 960 1 INV1S $T=982700 376440 1 0 $X=982700 $Y=371020
X404 5486 2 5442 1 INV1S $T=984560 426840 1 180 $X=983320 $Y=426460
X405 973 2 929 1 INV1S $T=990140 537720 0 180 $X=988900 $Y=532300
X406 5515 2 5510 1 INV1S $T=989520 487320 0 0 $X=989520 $Y=486940
X407 5479 2 980 1 INV1S $T=992000 406680 1 0 $X=992000 $Y=401260
X408 5460 2 5545 1 INV1S $T=993240 477240 1 0 $X=993240 $Y=471820
X409 5511 2 5486 1 INV1S $T=997580 426840 0 0 $X=997580 $Y=426460
X410 5555 2 5560 1 INV1S $T=997580 457080 0 0 $X=997580 $Y=456700
X411 5563 2 5571 1 INV1S $T=999440 416760 1 0 $X=999440 $Y=411340
X412 970 2 5440 1 INV1S $T=999440 487320 0 0 $X=999440 $Y=486940
X413 996 2 5594 1 INV1S $T=1003780 376440 1 0 $X=1003780 $Y=371020
X414 5486 2 5615 1 INV1S $T=1005020 426840 0 0 $X=1005020 $Y=426460
X415 5574 2 5603 1 INV1S $T=1005640 416760 0 0 $X=1005640 $Y=416380
X416 5467 2 5612 1 INV1S $T=1005640 507480 1 0 $X=1005640 $Y=502060
X417 5612 2 5570 1 INV1S $T=1006260 507480 0 0 $X=1006260 $Y=507100
X418 5500 2 5623 1 INV1S $T=1006880 477240 0 0 $X=1006880 $Y=476860
X419 5611 2 5644 1 INV1S $T=1011220 497400 1 0 $X=1011220 $Y=491980
X420 5614 2 5640 1 INV1S $T=1013700 396600 1 0 $X=1013700 $Y=391180
X421 5623 2 5658 1 INV1S $T=1020520 477240 1 180 $X=1019280 $Y=476860
X422 5669 2 5586 1 INV1S $T=1021140 467160 1 180 $X=1019900 $Y=466780
X423 5549 2 5676 1 INV1S $T=1020520 426840 0 0 $X=1020520 $Y=426460
X424 5670 2 5669 1 INV1S $T=1023000 467160 1 180 $X=1021760 $Y=466780
X425 5623 2 5687 1 INV1S $T=1024240 487320 1 0 $X=1024240 $Y=481900
X426 885 2 5727 1 INV1S $T=1031680 426840 0 0 $X=1031680 $Y=426460
X427 5753 2 5713 1 INV1S $T=1036020 396600 0 180 $X=1034780 $Y=391180
X428 5612 2 5762 1 INV1S $T=1039740 507480 0 0 $X=1039740 $Y=507100
X429 5594 2 5753 1 INV1S $T=1040360 396600 1 0 $X=1040360 $Y=391180
X430 5466 2 5800 1 INV1S $T=1045940 447000 1 0 $X=1045940 $Y=441580
X431 5753 2 5751 1 INV1S $T=1047180 396600 1 0 $X=1047180 $Y=391180
X432 5800 2 5768 1 INV1S $T=1048420 447000 1 0 $X=1048420 $Y=441580
X433 5676 2 5761 1 INV1S $T=1051520 426840 1 180 $X=1050280 $Y=426460
X434 1077 2 5853 1 INV1S $T=1058960 537720 1 0 $X=1058960 $Y=532300
X435 5676 2 5854 1 INV1S $T=1059580 426840 0 0 $X=1059580 $Y=426460
X436 5613 2 5884 1 INV1S $T=1066400 406680 0 0 $X=1066400 $Y=406300
X437 5800 2 5905 1 INV1S $T=1068880 436920 0 0 $X=1068880 $Y=436540
X438 5884 2 5896 1 INV1S $T=1075080 406680 0 0 $X=1075080 $Y=406300
X439 5988 2 1103 1 INV1S $T=1089340 507480 1 180 $X=1088100 $Y=507100
X440 1104 2 5988 1 INV1S $T=1088100 517560 1 0 $X=1088100 $Y=512140
X441 5988 2 5999 1 INV1S $T=1091820 507480 0 0 $X=1091820 $Y=507100
X442 5988 2 6003 1 INV1S $T=1093680 507480 1 0 $X=1093680 $Y=502060
X443 5680 2 6019 1 INV1S $T=1094920 416760 0 0 $X=1094920 $Y=416380
X444 5853 2 6080 1 INV1S $T=1107940 527640 0 0 $X=1107940 $Y=527260
X445 1076 2 5966 1 INV1S $T=1108560 527640 1 0 $X=1108560 $Y=522220
X446 1124 2 6099 1 INV1S $T=1115380 507480 1 180 $X=1114140 $Y=507100
X447 1124 2 1123 1 INV1S $T=1115380 426840 0 0 $X=1115380 $Y=426460
X448 1132 2 1135 1 INV1S $T=1127160 386520 1 0 $X=1127160 $Y=381100
X449 1135 2 6141 1 INV1S $T=1127780 406680 1 0 $X=1127780 $Y=401260
X450 1124 2 6027 1 INV1S $T=1127780 416760 1 0 $X=1127780 $Y=411340
X451 1219 1 2 1207 BUF1S $T=223200 457080 0 180 $X=220720 $Y=451660
X452 16 1 2 1208 BUF1S $T=223200 477240 1 180 $X=220720 $Y=476860
X453 1205 1 2 1209 BUF1S $T=223200 517560 1 180 $X=220720 $Y=517180
X454 14 1 2 5 BUF1S $T=223200 537720 0 180 $X=220720 $Y=532300
X455 12 1 2 1206 BUF1S $T=222580 416760 1 0 $X=222580 $Y=411340
X456 7 1 2 1230 BUF1S $T=222580 447000 1 0 $X=222580 $Y=441580
X457 1203 1 2 1235 BUF1S $T=223200 426840 1 0 $X=223200 $Y=421420
X458 1237 1 2 26 BUF1S $T=227540 376440 1 0 $X=227540 $Y=371020
X459 1207 1 2 21 BUF1S $T=227540 386520 1 0 $X=227540 $Y=381100
X460 1217 1 2 1264 BUF1S $T=227540 477240 0 0 $X=227540 $Y=476860
X461 1222 1 2 1289 BUF1S $T=232500 386520 0 0 $X=232500 $Y=386140
X462 1231 1 2 1280 BUF1S $T=233120 457080 1 0 $X=233120 $Y=451660
X463 1278 1 2 1297 BUF1S $T=234360 467160 0 0 $X=234360 $Y=466780
X464 1226 1 2 28 BUF1S $T=234980 376440 1 0 $X=234980 $Y=371020
X465 1240 1 2 1299 BUF1S $T=234980 436920 1 0 $X=234980 $Y=431500
X466 1309 1 2 1294 BUF1S $T=239320 426840 1 180 $X=236840 $Y=426460
X467 1219 1 2 1268 BUF1S $T=236840 447000 0 0 $X=236840 $Y=446620
X468 1241 1 2 1309 BUF1S $T=236840 457080 1 0 $X=236840 $Y=451660
X469 1280 1 2 1322 BUF1S $T=238700 406680 0 0 $X=238700 $Y=406300
X470 1293 1 2 1314 BUF1S $T=238700 487320 0 0 $X=238700 $Y=486940
X471 39 1 2 1250 BUF1S $T=242420 527640 1 180 $X=239940 $Y=527260
X472 1314 1 2 1320 BUF1S $T=241180 467160 0 0 $X=241180 $Y=466780
X473 1221 1 2 1346 BUF1S $T=243660 406680 0 0 $X=243660 $Y=406300
X474 1230 1 2 1353 BUF1S $T=243660 416760 0 0 $X=243660 $Y=416380
X475 43 1 2 41 BUF1S $T=246760 507480 0 180 $X=244280 $Y=502060
X476 1359 1 2 1338 BUF1S $T=248000 497400 1 180 $X=245520 $Y=497020
X477 47 1 2 1243 BUF1S $T=249240 527640 1 180 $X=246760 $Y=527260
X478 1385 1 2 1370 BUF1S $T=254820 497400 0 180 $X=252340 $Y=491980
X479 1235 1 2 1394 BUF1S $T=254200 386520 1 0 $X=254200 $Y=381100
X480 1392 1 2 1384 BUF1S $T=257920 497400 1 0 $X=257920 $Y=491980
X481 1395 1 2 1385 BUF1S $T=259780 527640 1 0 $X=259780 $Y=522220
X482 56 1 2 1420 BUF1S $T=264120 517560 1 180 $X=261640 $Y=517180
X483 60 1 2 48 BUF1S $T=262880 477240 0 0 $X=262880 $Y=476860
X484 64 1 2 46 BUF1S $T=267840 477240 1 180 $X=265360 $Y=476860
X485 63 1 2 1446 BUF1S $T=266600 517560 0 0 $X=266600 $Y=517180
X486 65 1 2 1453 BUF1S $T=274040 517560 0 180 $X=271560 $Y=512140
X487 1482 1 2 73 BUF1S $T=275900 376440 1 0 $X=275900 $Y=371020
X488 1505 1 2 68 BUF1S $T=280860 416760 1 0 $X=280860 $Y=411340
X489 79 1 2 1485 BUF1S $T=287060 527640 1 180 $X=284580 $Y=527260
X490 80 1 2 1486 BUF1S $T=287060 537720 0 180 $X=284580 $Y=532300
X491 1534 1 2 1482 BUF1S $T=288920 426840 0 180 $X=286440 $Y=421420
X492 1578 1 2 1505 BUF1S $T=293880 457080 1 180 $X=291400 $Y=456700
X493 1727 1 2 1745 BUF1S $T=312480 416760 0 0 $X=312480 $Y=416380
X494 1745 1 2 111 BUF1S $T=316820 376440 0 0 $X=316820 $Y=376060
X495 107 1 2 1776 BUF1S $T=316820 447000 0 0 $X=316820 $Y=446620
X496 1758 1 2 1785 BUF1S $T=318060 406680 0 0 $X=318060 $Y=406300
X497 1785 1 2 112 BUF1S $T=322400 376440 1 180 $X=319920 $Y=376060
X498 1795 1 2 1758 BUF1S $T=323020 467160 1 180 $X=320540 $Y=466780
X499 1578 1 2 1801 BUF1S $T=321160 467160 1 0 $X=321160 $Y=461740
X500 116 1 2 1787 BUF1S $T=323640 517560 1 0 $X=323640 $Y=512140
X501 1805 1 2 118 BUF1S $T=325500 386520 0 0 $X=325500 $Y=386140
X502 1837 1 2 1578 BUF1S $T=329840 487320 0 180 $X=327360 $Y=481900
X503 1787 1 2 1805 BUF1S $T=331700 436920 1 180 $X=329220 $Y=436540
X504 1840 1 2 1850 BUF1S $T=329840 426840 1 0 $X=329840 $Y=421420
X505 1801 1 2 1860 BUF1S $T=332320 426840 1 0 $X=332320 $Y=421420
X506 1860 1 2 122 BUF1S $T=336660 386520 0 180 $X=334180 $Y=381100
X507 1862 1 2 1866 BUF1S $T=334180 497400 0 0 $X=334180 $Y=497020
X508 125 1 2 1869 BUF1S $T=336660 497400 0 0 $X=336660 $Y=497020
X509 1853 1 2 126 BUF1S $T=341620 366360 1 180 $X=339140 $Y=365980
X510 1796 1 2 131 BUF1S $T=342240 386520 0 0 $X=342240 $Y=386140
X511 1967 1 2 1973 BUF1S $T=355880 467160 0 0 $X=355880 $Y=466780
X512 2046 1 2 1969 BUF1S $T=366420 457080 0 180 $X=363940 $Y=451660
X513 2062 1 2 1995 BUF1S $T=367660 477240 1 180 $X=365180 $Y=476860
X514 2091 1 2 2023 BUF1S $T=372620 457080 1 180 $X=370140 $Y=456700
X515 2145 1 2 2045 BUF1S $T=381300 426840 1 180 $X=378820 $Y=426460
X516 171 1 2 2153 BUF1S $T=384400 416760 1 0 $X=384400 $Y=411340
X517 2216 1 2 2092 BUF1S $T=391840 457080 0 180 $X=389360 $Y=451660
X518 2046 1 2 178 BUF1S $T=393080 416760 0 180 $X=390600 $Y=411340
X519 2091 1 2 174 BUF1S $T=391220 436920 1 0 $X=391220 $Y=431500
X520 184 1 2 1744 BUF1S $T=393700 527640 1 180 $X=391220 $Y=527260
X521 2225 1 2 187 BUF1S $T=393080 396600 0 0 $X=393080 $Y=396220
X522 2225 1 2 1967 BUF1S $T=398040 436920 1 180 $X=395560 $Y=436540
X523 2260 1 2 2037 BUF1S $T=398660 447000 1 180 $X=396180 $Y=446620
X524 2216 1 2 185 BUF1S $T=396800 426840 0 0 $X=396800 $Y=426460
X525 2267 1 2 2015 BUF1S $T=400520 457080 1 180 $X=398040 $Y=456700
X526 197 1 2 1980 BUF1S $T=402380 487320 0 180 $X=399900 $Y=481900
X527 2292 1 2 1972 BUF1S $T=404860 467160 1 180 $X=402380 $Y=466780
X528 2080 1 2 203 BUF1S $T=405480 527640 1 0 $X=405480 $Y=522220
X529 2347 1 2 212 BUF1S $T=412300 527640 1 0 $X=412300 $Y=522220
X530 2386 1 2 2080 BUF1S $T=420360 507480 1 0 $X=420360 $Y=502060
X531 2402 1 2 225 BUF1S $T=424700 386520 0 0 $X=424700 $Y=386140
X532 1862 1 2 230 BUF1S $T=427180 386520 0 0 $X=427180 $Y=386140
X533 2402 1 2 2409 BUF1S $T=427180 457080 0 0 $X=427180 $Y=456700
X534 2299 1 2 229 BUF1S $T=427800 447000 1 0 $X=427800 $Y=441580
X535 2374 1 2 232 BUF1S $T=430280 447000 1 0 $X=430280 $Y=441580
X536 2457 1 2 1795 BUF1S $T=433380 467160 1 180 $X=430900 $Y=466780
X537 2457 1 2 2408 BUF1S $T=433380 467160 0 0 $X=433380 $Y=466780
X538 2411 1 2 234 BUF1S $T=435240 447000 1 0 $X=435240 $Y=441580
X539 2399 1 2 2489 BUF1S $T=437100 477240 1 0 $X=437100 $Y=471820
X540 2375 1 2 235 BUF1S $T=440200 447000 0 180 $X=437720 $Y=441580
X541 2518 1 2 233 BUF1S $T=443300 416760 0 180 $X=440820 $Y=411340
X542 2457 1 2 249 BUF1S $T=445160 507480 0 180 $X=442680 $Y=502060
X543 2380 1 2 2507 BUF1S $T=445160 517560 1 0 $X=445160 $Y=512140
X544 244 1 2 2531 BUF1S $T=446400 386520 1 0 $X=446400 $Y=381100
X545 228 1 2 2574 BUF1S $T=449500 426840 0 0 $X=449500 $Y=426460
X546 2488 1 2 2570 BUF1S $T=449500 467160 0 0 $X=449500 $Y=466780
X547 256 1 2 2583 BUF1S $T=449500 497400 0 0 $X=449500 $Y=497020
X548 257 1 2 2576 BUF1S $T=450740 396600 1 0 $X=450740 $Y=391180
X549 2372 1 2 2564 BUF1S $T=450740 517560 0 0 $X=450740 $Y=517180
X550 266 1 2 2593 BUF1S $T=460040 386520 0 0 $X=460040 $Y=386140
X551 268 1 2 2637 BUF1S $T=462520 537720 1 0 $X=462520 $Y=532300
X552 1853 1 2 2646 BUF1S $T=463140 426840 1 0 $X=463140 $Y=421420
X553 1862 1 2 2664 BUF1S $T=465620 416760 1 0 $X=465620 $Y=411340
X554 2574 1 2 284 BUF1S $T=467480 396600 1 0 $X=467480 $Y=391180
X555 2583 1 2 2749 BUF1S $T=478640 507480 0 0 $X=478640 $Y=507100
X556 2555 1 2 297 BUF1S $T=480500 467160 1 0 $X=480500 $Y=461740
X557 304 1 2 271 BUF1S $T=485460 527640 0 180 $X=482980 $Y=522220
X558 2646 1 2 2735 BUF1S $T=485460 416760 1 0 $X=485460 $Y=411340
X559 2646 1 2 2783 BUF1S $T=485460 426840 0 0 $X=485460 $Y=426460
X560 312 1 2 2778 BUF1S $T=488560 537720 1 0 $X=488560 $Y=532300
X561 2813 1 2 320 BUF1S $T=492280 376440 0 0 $X=492280 $Y=376060
X562 2735 1 2 2813 BUF1S $T=492280 396600 0 0 $X=492280 $Y=396220
X563 2570 1 2 2825 BUF1S $T=492280 467160 0 0 $X=492280 $Y=466780
X564 2836 1 2 2809 BUF1S $T=496620 406680 1 180 $X=494140 $Y=406300
X565 2748 1 2 2811 BUF1S $T=494760 467160 0 0 $X=494760 $Y=466780
X566 2816 1 2 2834 BUF1S $T=498480 416760 0 180 $X=496000 $Y=411340
X567 2789 1 2 2855 BUF1S $T=496000 426840 0 0 $X=496000 $Y=426460
X568 2839 1 2 2857 BUF1S $T=496000 497400 0 0 $X=496000 $Y=497020
X569 2721 1 2 2860 BUF1S $T=497860 457080 1 0 $X=497860 $Y=451660
X570 2866 1 2 2723 BUF1S $T=500340 477240 1 180 $X=497860 $Y=476860
X571 2723 1 2 2867 BUF1S $T=497860 507480 1 0 $X=497860 $Y=502060
X572 2788 1 2 2870 BUF1S $T=499100 426840 1 0 $X=499100 $Y=421420
X573 2884 1 2 2869 BUF1S $T=503440 426840 1 180 $X=500960 $Y=426460
X574 2667 1 2 2839 BUF1S $T=500960 487320 0 0 $X=500960 $Y=486940
X575 2860 1 2 2884 BUF1S $T=501580 436920 0 0 $X=501580 $Y=436540
X576 2730 1 2 2895 BUF1S $T=502200 406680 1 0 $X=502200 $Y=401260
X577 327 1 2 2736 BUF1S $T=505300 497400 1 180 $X=502820 $Y=497020
X578 2837 1 2 2919 BUF1S $T=510260 436920 1 180 $X=507780 $Y=436540
X579 2895 1 2 2948 BUF1S $T=508400 406680 1 0 $X=508400 $Y=401260
X580 2847 1 2 2971 BUF1S $T=510880 477240 0 0 $X=510880 $Y=476860
X581 2884 1 2 2914 BUF1S $T=517080 426840 0 0 $X=517080 $Y=426460
X582 2880 1 2 3045 BUF1S $T=518940 416760 0 0 $X=518940 $Y=416380
X583 313 1 2 3042 BUF1S $T=519560 497400 1 0 $X=519560 $Y=491980
X584 2984 1 2 360 BUF1S $T=520180 376440 1 0 $X=520180 $Y=371020
X585 3049 1 2 3057 BUF1S $T=521420 527640 0 0 $X=521420 $Y=527260
X586 3045 1 2 2984 BUF1S $T=522660 386520 0 0 $X=522660 $Y=386140
X587 3092 1 2 3107 BUF1S $T=527620 497400 0 0 $X=527620 $Y=497020
X588 2919 1 2 3117 BUF1S $T=527620 517560 1 0 $X=527620 $Y=512140
X589 3008 1 2 3157 BUF1S $T=533200 396600 1 0 $X=533200 $Y=391180
X590 2836 1 2 3180 BUF1S $T=536920 406680 1 0 $X=536920 $Y=401260
X591 2855 1 2 3191 BUF1S $T=536920 436920 1 0 $X=536920 $Y=431500
X592 2986 1 2 3182 BUF1S $T=538780 406680 0 0 $X=538780 $Y=406300
X593 2847 1 2 3204 BUF1S $T=538780 477240 0 0 $X=538780 $Y=476860
X594 3048 1 2 3205 BUF1S $T=538780 497400 1 0 $X=538780 $Y=491980
X595 3054 1 2 3185 BUF1S $T=538780 517560 1 0 $X=538780 $Y=512140
X596 2749 1 2 387 BUF1S $T=538780 537720 1 0 $X=538780 $Y=532300
X597 3182 1 2 3213 BUF1S $T=544980 376440 1 180 $X=542500 $Y=376060
X598 365 1 2 3232 BUF1S $T=543120 527640 1 0 $X=543120 $Y=522220
X599 3204 1 2 3135 BUF1S $T=546220 497400 0 180 $X=543740 $Y=491980
X600 340 1 2 3238 BUF1S $T=545600 396600 0 0 $X=545600 $Y=396220
X601 2937 1 2 3253 BUF1S $T=547460 416760 0 0 $X=547460 $Y=416380
X602 3266 1 2 3134 BUF1S $T=551180 487320 0 180 $X=548700 $Y=481900
X603 341 1 2 3273 BUF1S $T=549940 416760 0 0 $X=549940 $Y=416380
X604 2948 1 2 399 BUF1S $T=551800 396600 1 0 $X=551800 $Y=391180
X605 3150 1 2 3247 BUF1S $T=551800 497400 0 0 $X=551800 $Y=497020
X606 2932 1 2 3298 BUF1S $T=552420 426840 0 0 $X=552420 $Y=426460
X607 3180 1 2 3296 BUF1S $T=556760 396600 0 0 $X=556760 $Y=396220
X608 3020 1 2 391 BUF1S $T=559240 497400 1 180 $X=556760 $Y=497020
X609 2921 1 2 3324 BUF1S $T=559860 426840 1 0 $X=559860 $Y=421420
X610 3104 1 2 401 BUF1S $T=562340 487320 0 180 $X=559860 $Y=481900
X611 3131 1 2 411 BUF1S $T=563580 396600 1 0 $X=563580 $Y=391180
X612 3273 1 2 412 BUF1S $T=563580 396600 0 0 $X=563580 $Y=396220
X613 3316 1 2 3360 BUF1S $T=563580 406680 1 0 $X=563580 $Y=401260
X614 413 1 2 3095 BUF1S $T=566680 517560 0 180 $X=564200 $Y=512140
X615 3360 1 2 419 BUF1S $T=573500 376440 0 180 $X=571020 $Y=371020
X616 3346 1 2 418 BUF1S $T=572260 366360 0 0 $X=572260 $Y=365980
X617 3408 1 2 3349 BUF1S $T=575360 487320 1 180 $X=572880 $Y=486940
X618 3413 1 2 3346 BUF1S $T=580320 406680 1 0 $X=580320 $Y=401260
X619 3572 1 2 3590 BUF1S $T=600780 457080 1 0 $X=600780 $Y=451660
X620 3408 1 2 3617 BUF1S $T=605740 517560 1 0 $X=605740 $Y=512140
X621 3630 1 2 3636 BUF1S $T=609460 467160 1 0 $X=609460 $Y=461740
X622 3608 1 2 3654 BUF1S $T=615660 467160 0 180 $X=613180 $Y=461740
X623 3680 1 2 461 BUF1S $T=621240 376440 1 180 $X=618760 $Y=376060
X624 3706 1 2 460 BUF1S $T=622480 396600 0 180 $X=620000 $Y=391180
X625 3823 1 2 3734 BUF1S $T=643560 386520 1 180 $X=641080 $Y=386140
X626 3831 1 2 3728 BUF1S $T=644180 386520 0 180 $X=641700 $Y=381100
X627 468 1 2 514 BUF1S $T=652240 366360 0 0 $X=652240 $Y=365980
X628 3917 1 2 3873 BUF1S $T=655960 406680 0 0 $X=655960 $Y=406300
X629 3995 1 2 523 BUF1S $T=670220 497400 1 180 $X=667740 $Y=497020
X630 531 1 2 4002 BUF1S $T=671460 527640 0 0 $X=671460 $Y=527260
X631 3948 1 2 3986 BUF1S $T=676420 487320 0 180 $X=673940 $Y=481900
X632 3986 1 2 4033 BUF1S $T=675180 477240 1 0 $X=675180 $Y=471820
X633 3972 1 2 3981 BUF1S $T=680760 517560 1 0 $X=680760 $Y=512140
X634 3972 1 2 4080 BUF1S $T=685100 517560 0 0 $X=685100 $Y=517180
X635 548 1 2 3963 BUF1S $T=690060 517560 1 180 $X=687580 $Y=517180
X636 4069 1 2 4056 BUF1S $T=699980 436920 0 180 $X=697500 $Y=431500
X637 4131 1 2 4138 BUF1S $T=701840 426840 1 180 $X=699360 $Y=426460
X638 4136 1 2 4069 BUF1S $T=704320 426840 1 180 $X=701840 $Y=426460
X639 564 1 2 4077 BUF1S $T=701840 507480 1 0 $X=701840 $Y=502060
X640 4136 1 2 4111 BUF1S $T=703700 396600 0 0 $X=703700 $Y=396220
X641 4179 1 2 4087 BUF1S $T=706180 457080 0 180 $X=703700 $Y=451660
X642 3981 1 2 4156 BUF1S $T=703700 497400 1 0 $X=703700 $Y=491980
X643 4173 1 2 4120 BUF1S $T=706180 517560 1 180 $X=703700 $Y=517180
X644 4188 1 2 4099 BUF1S $T=707420 477240 1 0 $X=707420 $Y=471820
X645 4197 1 2 4019 BUF1S $T=709900 497400 0 180 $X=707420 $Y=491980
X646 4210 1 2 4105 BUF1S $T=713620 447000 0 180 $X=711140 $Y=441580
X647 4192 1 2 4215 BUF1S $T=712380 376440 0 0 $X=712380 $Y=376060
X648 4205 1 2 4119 BUF1S $T=715480 467160 1 180 $X=713000 $Y=466780
X649 4220 1 2 4036 BUF1S $T=716100 457080 1 180 $X=713620 $Y=456700
X650 4231 1 2 4118 BUF1S $T=716720 416760 1 180 $X=714240 $Y=416380
X651 4136 1 2 4223 BUF1S $T=714240 426840 1 0 $X=714240 $Y=421420
X652 582 1 2 4053 BUF1S $T=716720 527640 1 180 $X=714240 $Y=527260
X653 4136 1 2 572 BUF1S $T=716100 386520 0 0 $X=716100 $Y=386140
X654 4239 1 2 4146 BUF1S $T=720440 406680 0 180 $X=717960 $Y=401260
X655 4080 1 2 4226 BUF1S $T=719820 517560 0 0 $X=719820 $Y=517180
X656 4268 1 2 4089 BUF1S $T=724160 426840 1 180 $X=721680 $Y=426460
X657 4276 1 2 3967 BUF1S $T=726020 517560 1 180 $X=723540 $Y=517180
X658 575 1 2 4214 BUF1S $T=728500 386520 1 0 $X=728500 $Y=381100
X659 4322 1 2 4172 BUF1S $T=738420 376440 1 180 $X=735940 $Y=376060
X660 4324 1 2 4022 BUF1S $T=740280 457080 1 180 $X=737800 $Y=456700
X661 4223 1 2 4323 BUF1S $T=739040 406680 1 0 $X=739040 $Y=401260
X662 4303 1 2 4237 BUF1S $T=742140 457080 0 180 $X=739660 $Y=451660
X663 607 1 2 4353 BUF1S $T=740900 537720 1 0 $X=740900 $Y=532300
X664 4315 1 2 4359 BUF1S $T=742760 406680 1 0 $X=742760 $Y=401260
X665 4215 1 2 615 BUF1S $T=744620 376440 0 0 $X=744620 $Y=376060
X666 618 1 2 4206 BUF1S $T=748960 386520 0 180 $X=746480 $Y=381100
X667 564 1 2 4382 BUF1S $T=746480 517560 0 0 $X=746480 $Y=517180
X668 4324 1 2 4385 BUF1S $T=747100 447000 1 0 $X=747100 $Y=441580
X669 616 1 2 4388 BUF1S $T=748340 457080 1 0 $X=748340 $Y=451660
X670 4404 1 2 4338 BUF1S $T=750820 477240 0 180 $X=748340 $Y=471820
X671 4231 1 2 4401 BUF1S $T=750200 406680 0 0 $X=750200 $Y=406300
X672 4197 1 2 4400 BUF1S $T=750200 497400 1 0 $X=750200 $Y=491980
X673 4322 1 2 627 BUF1S $T=752060 376440 0 0 $X=752060 $Y=376060
X674 4315 1 2 4339 BUF1S $T=752060 436920 0 0 $X=752060 $Y=436540
X675 4173 1 2 629 BUF1S $T=753300 527640 0 0 $X=753300 $Y=527260
X676 4220 1 2 4415 BUF1S $T=753920 447000 1 0 $X=753920 $Y=441580
X677 4268 1 2 4430 BUF1S $T=757020 426840 1 0 $X=757020 $Y=421420
X678 4210 1 2 4444 BUF1S $T=757020 426840 0 0 $X=757020 $Y=426460
X679 4205 1 2 4426 BUF1S $T=757020 467160 0 0 $X=757020 $Y=466780
X680 4239 1 2 4356 BUF1S $T=758260 396600 0 0 $X=758260 $Y=396220
X681 4456 1 2 4159 BUF1S $T=763840 406680 0 180 $X=761360 $Y=401260
X682 4404 1 2 4481 BUF1S $T=767560 457080 0 0 $X=767560 $Y=456700
X683 4483 1 2 614 BUF1S $T=771280 527640 1 180 $X=768800 $Y=527260
X684 4518 1 2 4414 BUF1S $T=773140 396600 0 180 $X=770660 $Y=391180
X685 4276 1 2 4513 BUF1S $T=771900 507480 1 0 $X=771900 $Y=502060
X686 3995 1 2 4524 BUF1S $T=774380 497400 0 0 $X=774380 $Y=497020
X687 613 1 2 4496 BUF1S $T=775620 527640 0 0 $X=775620 $Y=527260
X688 4481 1 2 4539 BUF1S $T=792360 447000 0 0 $X=792360 $Y=446620
X689 662 1 2 4464 BUF1S $T=796700 507480 1 180 $X=794220 $Y=507100
X690 651 1 2 4635 BUF1S $T=799800 507480 1 0 $X=799800 $Y=502060
X691 4570 1 2 4591 BUF1S $T=801660 416760 0 0 $X=801660 $Y=416380
X692 4423 1 2 4610 BUF1S $T=812200 477240 0 0 $X=812200 $Y=476860
X693 4704 1 2 4626 BUF1S $T=816540 447000 1 180 $X=814060 $Y=446620
X694 591 1 2 4742 BUF1S $T=822740 426840 0 0 $X=822740 $Y=426460
X695 4717 1 2 4670 BUF1S $T=825840 406680 0 180 $X=823360 $Y=401260
X696 4642 1 2 4719 BUF1S $T=824600 517560 0 0 $X=824600 $Y=517180
X697 4754 1 2 4728 BUF1S $T=828940 436920 0 180 $X=826460 $Y=431500
X698 4704 1 2 4751 BUF1S $T=828320 447000 1 0 $X=828320 $Y=441580
X699 4752 1 2 4739 BUF1S $T=830800 467160 0 180 $X=828320 $Y=461740
X700 698 1 2 4642 BUF1S $T=833900 527640 1 180 $X=831420 $Y=527260
X701 4717 1 2 4743 BUF1S $T=832040 416760 0 0 $X=832040 $Y=416380
X702 4722 1 2 4768 BUF1S $T=832660 487320 0 0 $X=832660 $Y=486940
X703 4779 1 2 4725 BUF1S $T=837620 416760 0 180 $X=835140 $Y=411340
X704 4751 1 2 4722 BUF1S $T=835140 467160 1 0 $X=835140 $Y=461740
X705 4779 1 2 4805 BUF1S $T=838240 416760 1 0 $X=838240 $Y=411340
X706 4781 1 2 4776 BUF1S $T=841340 487320 1 180 $X=838860 $Y=486940
X707 4743 1 2 4756 BUF1S $T=845060 396600 0 180 $X=842580 $Y=391180
X708 705 1 2 4812 BUF1S $T=842580 527640 1 0 $X=842580 $Y=522220
X709 4754 1 2 4830 BUF1S $T=844440 426840 0 0 $X=844440 $Y=426460
X710 4743 1 2 4845 BUF1S $T=847540 416760 1 0 $X=847540 $Y=411340
X711 4841 1 2 4820 BUF1S $T=850020 497400 1 180 $X=847540 $Y=497020
X712 4597 1 2 745 BUF1S $T=851260 406680 1 0 $X=851260 $Y=401260
X713 4751 1 2 4863 BUF1S $T=851260 447000 0 0 $X=851260 $Y=446620
X714 4768 1 2 4787 BUF1S $T=856840 507480 0 180 $X=854360 $Y=502060
X715 757 1 2 735 BUF1S $T=856840 527640 1 180 $X=854360 $Y=527260
X716 4865 1 2 4858 BUF1S $T=857460 477240 0 180 $X=854980 $Y=471820
X717 619 1 2 4895 BUF1S $T=856840 467160 0 0 $X=856840 $Y=466780
X718 4926 1 2 4876 BUF1S $T=862420 477240 1 180 $X=859940 $Y=476860
X719 769 1 2 767 BUF1S $T=863040 366360 1 180 $X=860560 $Y=365980
X720 4915 1 2 4898 BUF1S $T=864900 517560 1 180 $X=862420 $Y=517180
X721 4928 1 2 4883 BUF1S $T=863660 406680 0 0 $X=863660 $Y=406300
X722 602 1 2 4940 BUF1S $T=863660 426840 1 0 $X=863660 $Y=421420
X723 4941 1 2 4872 BUF1S $T=866140 436920 0 180 $X=863660 $Y=431500
X724 4768 1 2 4935 BUF1S $T=863660 477240 0 0 $X=863660 $Y=476860
X725 4941 1 2 4875 BUF1S $T=871720 376440 1 180 $X=869240 $Y=376060
X726 4958 1 2 4922 BUF1S $T=872960 406680 0 180 $X=870480 $Y=401260
X727 4863 1 2 4989 BUF1S $T=874200 447000 0 0 $X=874200 $Y=446620
X728 4845 1 2 4893 BUF1S $T=881640 416760 0 0 $X=881640 $Y=416380
X729 4935 1 2 5023 BUF1S $T=881640 477240 1 0 $X=881640 $Y=471820
X730 4739 1 2 5027 BUF1S $T=884740 477240 0 0 $X=884740 $Y=476860
X731 5014 1 2 808 BUF1S $T=885360 396600 1 0 $X=885360 $Y=391180
X732 4971 1 2 5048 BUF1S $T=886600 477240 1 0 $X=886600 $Y=471820
X733 5033 1 2 800 BUF1S $T=889700 386520 1 180 $X=887220 $Y=386140
X734 5045 1 2 5037 BUF1S $T=887840 527640 0 0 $X=887840 $Y=527260
X735 809 1 2 769 BUF1S $T=894660 366360 1 180 $X=892180 $Y=365980
X736 757 1 2 5091 BUF1S $T=896520 406680 1 0 $X=896520 $Y=401260
X737 4964 1 2 5104 BUF1S $T=899000 477240 1 0 $X=899000 $Y=471820
X738 4893 1 2 5081 BUF1S $T=905200 406680 1 180 $X=902720 $Y=406300
X739 4883 1 2 5122 BUF1S $T=904580 396600 1 0 $X=904580 $Y=391180
X740 5027 1 2 5138 BUF1S $T=904580 467160 1 0 $X=904580 $Y=461740
X741 4941 1 2 5154 BUF1S $T=905820 436920 1 0 $X=905820 $Y=431500
X742 5092 1 2 5127 BUF1S $T=907680 457080 0 0 $X=907680 $Y=456700
X743 4922 1 2 5212 BUF1S $T=916360 406680 1 0 $X=916360 $Y=401260
X744 4841 1 2 5192 BUF1S $T=916980 507480 1 0 $X=916980 $Y=502060
X745 790 1 2 5098 BUF1S $T=916980 527640 0 0 $X=916980 $Y=527260
X746 830 1 2 819 BUF1S $T=918840 467160 1 0 $X=918840 $Y=461740
X747 4830 1 2 5222 BUF1S $T=922560 396600 0 0 $X=922560 $Y=396220
X748 4891 1 2 5242 BUF1S $T=923800 376440 1 0 $X=923800 $Y=371020
X749 5192 1 2 5241 BUF1S $T=923800 457080 0 0 $X=923800 $Y=456700
X750 4805 1 2 5235 BUF1S $T=924420 396600 1 0 $X=924420 $Y=391180
X751 821 1 2 5249 BUF1S $T=925660 507480 0 0 $X=925660 $Y=507100
X752 4951 1 2 850 BUF1S $T=926280 376440 1 0 $X=926280 $Y=371020
X753 5126 1 2 5265 BUF1S $T=927520 477240 1 0 $X=927520 $Y=471820
X754 5266 1 2 5158 BUF1S $T=931860 436920 0 180 $X=929380 $Y=431500
X755 4876 1 2 5259 BUF1S $T=929380 507480 1 0 $X=929380 $Y=502060
X756 830 1 2 5219 BUF1S $T=933100 497400 0 180 $X=930620 $Y=491980
X757 757 1 2 5272 BUF1S $T=931240 406680 0 0 $X=931240 $Y=406300
X758 5143 1 2 5286 BUF1S $T=931860 386520 0 0 $X=931860 $Y=386140
X759 864 1 2 5133 BUF1S $T=934340 477240 1 0 $X=934340 $Y=471820
X760 5122 1 2 5292 BUF1S $T=936820 416760 1 0 $X=936820 $Y=411340
X761 4915 1 2 5321 BUF1S $T=941780 517560 1 0 $X=941780 $Y=512140
X762 5328 1 2 5236 BUF1S $T=946120 416760 0 180 $X=943640 $Y=411340
X763 5048 1 2 5338 BUF1S $T=943640 477240 1 0 $X=943640 $Y=471820
X764 871 1 2 5344 BUF1S $T=944260 487320 0 0 $X=944260 $Y=486940
X765 5104 1 2 5332 BUF1S $T=950460 477240 1 0 $X=950460 $Y=471820
X766 5254 1 2 5285 BUF1S $T=952940 507480 1 180 $X=950460 $Y=507100
X767 5261 1 2 5376 BUF1S $T=954180 477240 1 0 $X=954180 $Y=471820
X768 5376 1 2 5254 BUF1S $T=958520 477240 1 180 $X=956040 $Y=476860
X769 5289 1 2 5388 BUF1S $T=956040 487320 0 0 $X=956040 $Y=486940
X770 5364 1 2 5328 BUF1S $T=959760 416760 1 0 $X=959760 $Y=411340
X771 5321 1 2 5403 BUF1S $T=959760 477240 0 0 $X=959760 $Y=476860
X772 5259 1 2 5402 BUF1S $T=959760 507480 1 0 $X=959760 $Y=502060
X773 5212 1 2 5369 BUF1S $T=960380 406680 0 0 $X=960380 $Y=406300
X774 5364 1 2 5266 BUF1S $T=965340 426840 0 180 $X=962860 $Y=421420
X775 5376 1 2 5408 BUF1S $T=965340 477240 1 0 $X=965340 $Y=471820
X776 5381 1 2 917 BUF1S $T=969060 366360 1 180 $X=966580 $Y=365980
X777 5379 1 2 5381 BUF1S $T=966580 386520 1 0 $X=966580 $Y=381100
X778 5328 1 2 5379 BUF1S $T=969060 406680 1 180 $X=966580 $Y=406300
X779 5364 1 2 5429 BUF1S $T=966580 426840 1 0 $X=966580 $Y=421420
X780 5381 1 2 926 BUF1S $T=968440 376440 1 0 $X=968440 $Y=371020
X781 5429 1 2 5456 BUF1S $T=978980 436920 1 0 $X=978980 $Y=431500
X782 5510 1 2 5454 BUF1S $T=988900 507480 1 180 $X=986420 $Y=507100
X783 975 1 2 5538 BUF1S $T=990140 537720 1 0 $X=990140 $Y=532300
X784 5444 1 2 5549 BUF1S $T=991380 426840 0 0 $X=991380 $Y=426460
X785 5328 1 2 5547 BUF1S $T=993240 406680 1 0 $X=993240 $Y=401260
X786 5519 1 2 978 BUF1S $T=995100 457080 0 0 $X=995100 $Y=456700
X787 5571 1 2 5475 BUF1S $T=1001300 406680 1 180 $X=998820 $Y=406300
X788 5545 1 2 5556 BUF1S $T=999440 487320 1 0 $X=999440 $Y=481900
X789 5568 1 2 5592 BUF1S $T=1000060 467160 0 0 $X=1000060 $Y=466780
X790 5573 1 2 5481 BUF1S $T=1005020 416760 0 180 $X=1002540 $Y=411340
X791 5599 1 2 957 BUF1S $T=1005020 507480 1 180 $X=1002540 $Y=507100
X792 5603 1 2 5468 BUF1S $T=1006260 396600 1 180 $X=1003780 $Y=396220
X793 5510 1 2 5642 BUF1S $T=1006880 507480 1 0 $X=1006880 $Y=502060
X794 5429 1 2 5628 BUF1S $T=1011840 426840 0 0 $X=1011840 $Y=426460
X795 5556 1 2 5651 BUF1S $T=1013080 477240 0 0 $X=1013080 $Y=476860
X796 5640 1 2 1020 BUF1S $T=1018040 376440 0 0 $X=1018040 $Y=376060
X797 5674 1 2 5577 BUF1S $T=1021140 527640 1 180 $X=1018660 $Y=527260
X798 5596 1 2 1025 BUF1S $T=1020520 376440 1 0 $X=1020520 $Y=371020
X799 5457 1 2 5681 BUF1S $T=1021760 447000 1 0 $X=1021760 $Y=441580
X800 5577 1 2 5690 BUF1S $T=1021760 507480 0 0 $X=1021760 $Y=507100
X801 5560 1 2 5699 BUF1S $T=1027340 467160 0 0 $X=1027340 $Y=466780
X802 942 1 2 1042 BUF1S $T=1030440 376440 1 0 $X=1030440 $Y=371020
X803 5727 1 2 5748 BUF1S $T=1037880 447000 1 0 $X=1037880 $Y=441580
X804 1057 1 2 5674 BUF1S $T=1040360 527640 0 180 $X=1037880 $Y=522220
X805 5527 1 2 5771 BUF1S $T=1038500 467160 0 0 $X=1038500 $Y=466780
X806 1057 1 2 5788 BUF1S $T=1043460 527640 1 0 $X=1043460 $Y=522220
X807 1058 1 2 5765 BUF1S $T=1044080 527640 0 0 $X=1044080 $Y=527260
X808 5571 1 2 5789 BUF1S $T=1044700 406680 1 0 $X=1044700 $Y=401260
X809 5603 1 2 5790 BUF1S $T=1044700 406680 0 0 $X=1044700 $Y=406300
X810 980 1 2 1061 BUF1S $T=1047180 366360 0 0 $X=1047180 $Y=365980
X811 5615 1 2 5810 BUF1S $T=1048420 426840 1 0 $X=1048420 $Y=421420
X812 5519 1 2 5787 BUF1S $T=1049040 447000 0 0 $X=1049040 $Y=446620
X813 5727 1 2 5723 BUF1S $T=1054000 426840 1 180 $X=1051520 $Y=426460
X814 5687 1 2 5836 BUF1S $T=1054620 517560 1 0 $X=1054620 $Y=512140
X815 5642 1 2 5842 BUF1S $T=1055860 497400 1 0 $X=1055860 $Y=491980
X816 5644 1 2 5852 BUF1S $T=1057720 517560 0 0 $X=1057720 $Y=517180
X817 5723 1 2 5834 BUF1S $T=1061440 406680 1 180 $X=1058960 $Y=406300
X818 5762 1 2 5858 BUF1S $T=1058960 507480 0 0 $X=1058960 $Y=507100
X819 1080 1 2 5859 BUF1S $T=1060200 527640 1 0 $X=1060200 $Y=522220
X820 5596 1 2 1083 BUF1S $T=1062060 376440 0 0 $X=1062060 $Y=376060
X821 5727 1 2 5848 BUF1S $T=1064540 436920 0 0 $X=1064540 $Y=436540
X822 5681 1 2 5880 BUF1S $T=1064540 447000 0 0 $X=1064540 $Y=446620
X823 5699 1 2 5881 BUF1S $T=1064540 477240 1 0 $X=1064540 $Y=471820
X824 5771 1 2 5900 BUF1S $T=1067020 477240 1 0 $X=1067020 $Y=471820
X825 5410 1 2 5907 BUF1S $T=1067020 527640 1 0 $X=1067020 $Y=522220
X826 5848 1 2 5845 BUF1S $T=1070740 457080 0 180 $X=1068260 $Y=451660
X827 5834 1 2 5913 BUF1S $T=1069500 406680 1 0 $X=1069500 $Y=401260
X828 5788 1 2 5807 BUF1S $T=1070740 517560 1 0 $X=1070740 $Y=512140
X829 5848 1 2 5950 BUF1S $T=1084380 436920 0 180 $X=1081900 $Y=431500
X830 5845 1 2 5951 BUF1S $T=1091200 467160 0 180 $X=1088720 $Y=461740
X831 5913 1 2 5957 BUF1S $T=1101740 386520 1 0 $X=1101740 $Y=381100
X832 5950 1 2 6011 BUF1S $T=1103600 447000 1 0 $X=1103600 $Y=441580
X833 5950 1 2 5990 BUF1S $T=1104840 426840 0 0 $X=1104840 $Y=426460
X834 5990 1 2 6033 BUF1S $T=1107320 426840 0 0 $X=1107320 $Y=426460
X835 6011 1 2 6125 BUF1S $T=1114140 467160 0 0 $X=1114140 $Y=466780
X836 6033 1 2 1126 BUF1S $T=1120340 416760 1 0 $X=1120340 $Y=411340
X837 1121 1 2 6138 BUF1S $T=1124680 527640 1 0 $X=1124680 $Y=522220
X838 6141 1 2 1134 BUF1S $T=1129020 447000 1 180 $X=1126540 $Y=446620
X839 1234 1 2 1210 DELB $T=235600 527640 1 0 $X=235600 $Y=522220
X840 2675 1 2 2682 DELB $T=468100 487320 1 0 $X=468100 $Y=481900
X841 2726 1 2 2754 DELB $T=477400 457080 0 0 $X=477400 $Y=456700
X842 2784 1 2 2782 DELB $T=487320 457080 0 0 $X=487320 $Y=456700
X843 2792 1 2 2822 DELB $T=489180 426840 1 0 $X=489180 $Y=421420
X844 2796 1 2 2790 DELB $T=489180 517560 1 0 $X=489180 $Y=512140
X845 2824 1 2 2845 DELB $T=494140 457080 0 0 $X=494140 $Y=456700
X846 2858 1 2 2886 DELB $T=498480 517560 1 0 $X=498480 $Y=512140
X847 2864 1 2 2872 DELB $T=501580 467160 1 0 $X=501580 $Y=461740
X848 3667 1 2 3693 DELB $T=613800 487320 1 0 $X=613800 $Y=481900
X849 471 1 2 478 DELB $T=626200 467160 1 0 $X=626200 $Y=461740
X850 3874 1 2 3899 DELB $T=648520 497400 0 0 $X=648520 $Y=497020
X851 3893 1 2 3924 DELB $T=651620 527640 0 0 $X=651620 $Y=527260
X852 522 1 2 530 DELB $T=665880 406680 1 0 $X=665880 $Y=401260
X853 526 1 2 534 DELB $T=668980 416760 1 0 $X=668980 $Y=411340
X854 4004 1 2 4034 DELB $T=672700 487320 0 0 $X=672700 $Y=486940
X855 4062 1 2 4091 DELB $T=688820 477240 1 0 $X=688820 $Y=471820
X856 4104 1 2 4114 DELB $T=690680 436920 0 0 $X=690680 $Y=436540
X857 4054 1 2 558 DELB $T=691920 527640 0 0 $X=691920 $Y=527260
X858 4096 1 2 4128 DELB $T=695020 477240 0 0 $X=695020 $Y=476860
X859 4109 1 2 4171 DELB $T=698740 527640 0 0 $X=698740 $Y=527260
X860 4160 1 2 4187 DELB $T=706180 436920 0 0 $X=706180 $Y=436540
X861 4191 1 2 4196 DELB $T=707420 386520 1 0 $X=707420 $Y=381100
X862 4212 1 2 4213 DELB $T=713000 436920 0 0 $X=713000 $Y=436540
X863 4217 1 2 4218 DELB $T=714860 477240 0 0 $X=714860 $Y=476860
X864 4247 1 2 4274 DELB $T=721060 477240 1 0 $X=721060 $Y=471820
X865 4235 1 2 4249 DELB $T=721680 507480 0 0 $X=721680 $Y=507100
X866 4222 1 2 4230 DELB $T=723540 416760 0 0 $X=723540 $Y=416380
X867 4293 1 2 4321 DELB $T=730360 507480 0 0 $X=730360 $Y=507100
X868 4314 1 2 4335 DELB $T=733460 416760 0 0 $X=733460 $Y=416380
X869 4260 1 2 4308 DELB $T=737180 477240 1 0 $X=737180 $Y=471820
X870 4302 1 2 4341 DELB $T=739660 376440 1 0 $X=739660 $Y=371020
X871 4352 1 2 4358 DELB $T=742760 416760 0 0 $X=742760 $Y=416380
X872 4374 1 2 4376 DELB $T=747100 376440 0 0 $X=747100 $Y=376060
X873 4326 1 2 4331 DELB $T=747100 467160 1 0 $X=747100 $Y=461740
X874 4329 1 2 4343 DELB $T=747100 507480 0 0 $X=747100 $Y=507100
X875 4325 1 2 4381 DELB $T=748960 487320 1 0 $X=748960 $Y=481900
X876 4369 1 2 4405 DELB $T=753300 396600 0 0 $X=753300 $Y=396220
X877 4395 1 2 4393 DELB $T=755780 457080 1 0 $X=755780 $Y=451660
X878 4422 1 2 4439 DELB $T=757020 416760 1 0 $X=757020 $Y=411340
X879 4420 1 2 4424 DELB $T=757020 487320 1 0 $X=757020 $Y=481900
X880 4367 1 2 4411 DELB $T=759500 376440 0 0 $X=759500 $Y=376060
X881 4364 1 2 4357 DELB $T=759500 426840 1 0 $X=759500 $Y=421420
X882 4440 1 2 4463 DELB $T=761360 457080 1 0 $X=761360 $Y=451660
X883 4403 1 2 4452 DELB $T=764460 386520 1 0 $X=764460 $Y=381100
X884 4471 1 2 4478 DELB $T=767560 426840 1 0 $X=767560 $Y=421420
X885 4479 1 2 4509 DELB $T=768800 517560 0 0 $X=768800 $Y=517180
X886 4484 1 2 4491 DELB $T=770040 386520 1 0 $X=770040 $Y=381100
X887 4480 1 2 4492 DELB $T=771280 447000 0 0 $X=771280 $Y=446620
X888 4506 1 2 4529 DELB $T=773140 416760 0 0 $X=773140 $Y=416380
X889 4519 1 2 4538 DELB $T=775000 396600 0 0 $X=775000 $Y=396220
X890 4505 1 2 4487 DELB $T=775000 517560 1 0 $X=775000 $Y=512140
X891 4460 1 2 4474 DELB $T=776860 487320 0 0 $X=776860 $Y=486940
X892 4502 1 2 4540 DELB $T=780580 447000 0 0 $X=780580 $Y=446620
X893 4489 1 2 4534 DELB $T=782440 416760 0 0 $X=782440 $Y=416380
X894 4568 1 2 4574 DELB $T=789260 416760 0 0 $X=789260 $Y=416380
X895 4580 1 2 4605 DELB $T=792360 436920 0 0 $X=792360 $Y=436540
X896 4533 1 2 4541 DELB $T=792360 467160 1 0 $X=792360 $Y=461740
X897 4592 1 2 4598 DELB $T=794840 447000 0 0 $X=794840 $Y=446620
X898 4583 1 2 4596 DELB $T=795460 416760 1 0 $X=795460 $Y=411340
X899 4620 1 2 4625 DELB $T=801040 467160 1 0 $X=801040 $Y=461740
X900 4637 1 2 4662 DELB $T=802900 416760 1 0 $X=802900 $Y=411340
X901 4644 1 2 4638 DELB $T=804140 447000 0 0 $X=804140 $Y=446620
X902 4672 1 2 4676 DELB $T=810340 426840 1 0 $X=810340 $Y=421420
X903 4646 1 2 4654 DELB $T=814060 406680 0 0 $X=814060 $Y=406300
X904 4659 1 2 4658 DELB $T=816540 447000 0 0 $X=816540 $Y=446620
X905 4694 1 2 4702 DELB $T=817160 517560 0 0 $X=817160 $Y=517180
X906 4653 1 2 4693 DELB $T=822120 517560 1 0 $X=822120 $Y=512140
X907 4579 1 2 4588 DELB $T=825220 457080 1 0 $X=825220 $Y=451660
X908 4730 1 2 4741 DELB $T=826460 386520 1 0 $X=826460 $Y=381100
X909 4733 1 2 4753 DELB $T=830180 477240 0 0 $X=830180 $Y=476860
X910 4772 1 2 4764 DELB $T=834520 416760 0 0 $X=834520 $Y=416380
X911 4770 1 2 4775 DELB $T=835760 386520 1 0 $X=835760 $Y=381100
X912 4729 1 2 4782 DELB $T=835760 527640 1 0 $X=835760 $Y=522220
X913 4801 1 2 4819 DELB $T=838860 477240 1 0 $X=838860 $Y=471820
X914 4808 1 2 4832 DELB $T=842580 416760 1 0 $X=842580 $Y=411340
X915 4817 1 2 4833 DELB $T=842580 447000 0 0 $X=842580 $Y=446620
X916 4800 1 2 4821 DELB $T=843820 487320 1 0 $X=843820 $Y=481900
X917 737 1 2 4831 DELB $T=846920 376440 1 0 $X=846920 $Y=371020
X918 4834 1 2 4838 DELB $T=848780 396600 1 0 $X=848780 $Y=391180
X919 4763 1 2 4856 DELB $T=851260 457080 0 0 $X=851260 $Y=456700
X920 4843 1 2 4884 DELB $T=853740 436920 1 0 $X=853740 $Y=431500
X921 4889 1 2 4878 DELB $T=862420 517560 1 0 $X=862420 $Y=512140
X922 4908 1 2 4938 DELB $T=864280 376440 0 0 $X=864280 $Y=376060
X923 4946 1 2 4966 DELB $T=867380 366360 0 0 $X=867380 $Y=365980
X924 4950 1 2 4980 DELB $T=869860 426840 1 0 $X=869860 $Y=421420
X925 4953 1 2 4961 DELB $T=871100 517560 1 0 $X=871100 $Y=512140
X926 4987 1 2 5006 DELB $T=875440 426840 0 0 $X=875440 $Y=426460
X927 4984 1 2 5018 DELB $T=881020 376440 0 0 $X=881020 $Y=376060
X928 5042 1 2 5063 DELB $T=889080 477240 0 0 $X=889080 $Y=476860
X929 5071 1 2 5072 DELB $T=892800 396600 1 0 $X=892800 $Y=391180
X930 4998 1 2 5041 DELB $T=892800 477240 1 0 $X=892800 $Y=471820
X931 5085 1 2 5077 DELB $T=896520 507480 1 0 $X=896520 $Y=502060
X932 5119 1 2 5144 DELB $T=902720 477240 1 0 $X=902720 $Y=471820
X933 5093 1 2 5117 DELB $T=903960 396600 0 0 $X=903960 $Y=396220
X934 5111 1 2 5148 DELB $T=907680 416760 0 0 $X=907680 $Y=416380
X935 5112 1 2 5166 DELB $T=912020 396600 1 0 $X=912020 $Y=391180
X936 5174 1 2 5194 DELB $T=912020 507480 0 0 $X=912020 $Y=507100
X937 5141 1 2 5175 DELB $T=915740 517560 1 0 $X=915740 $Y=512140
X938 5186 1 2 5191 DELB $T=916360 416760 0 0 $X=916360 $Y=416380
X939 5171 1 2 5189 DELB $T=923180 457080 1 0 $X=923180 $Y=451660
X940 5230 1 2 5232 DELB $T=923800 426840 1 0 $X=923800 $Y=421420
X941 5237 1 2 5238 DELB $T=925040 487320 1 0 $X=925040 $Y=481900
X942 5198 1 2 5239 DELB $T=926900 396600 1 0 $X=926900 $Y=391180
X943 5244 1 2 5255 DELB $T=927520 517560 0 0 $X=927520 $Y=517180
X944 5270 1 2 5290 DELB $T=932480 487320 1 0 $X=932480 $Y=481900
X945 5264 1 2 5279 DELB $T=933720 396600 1 0 $X=933720 $Y=391180
X946 870 1 2 879 DELB $T=937440 366360 0 0 $X=937440 $Y=365980
X947 5310 1 2 5312 DELB $T=940540 426840 0 0 $X=940540 $Y=426460
X948 5314 1 2 5318 DELB $T=941780 467160 0 0 $X=941780 $Y=466780
X949 876 1 2 5322 DELB $T=947360 376440 1 0 $X=947360 $Y=371020
X950 5102 1 2 5109 DELB $T=947360 396600 0 0 $X=947360 $Y=396220
X951 5311 1 2 5300 DELB $T=947980 426840 0 0 $X=947980 $Y=426460
X952 5274 1 2 5304 DELB $T=951080 457080 1 0 $X=951080 $Y=451660
X953 5343 1 2 5356 DELB $T=951700 497400 0 0 $X=951700 $Y=497020
X954 5339 1 2 5360 DELB $T=952320 527640 0 0 $X=952320 $Y=527260
X955 5335 1 2 5363 DELB $T=953560 396600 0 0 $X=953560 $Y=396220
X956 5361 1 2 5371 DELB $T=955420 436920 1 0 $X=955420 $Y=431500
X957 5110 1 2 5120 DELB $T=955420 457080 0 0 $X=955420 $Y=456700
X958 5340 1 2 5404 DELB $T=957280 497400 0 0 $X=957280 $Y=497020
X959 5359 1 2 5366 DELB $T=957900 386520 1 0 $X=957900 $Y=381100
X960 5365 1 2 5368 DELB $T=957900 467160 1 0 $X=957900 $Y=461740
X961 5392 1 2 5421 DELB $T=965960 396600 1 0 $X=965960 $Y=391180
X962 5374 1 2 5424 DELB $T=967200 507480 0 0 $X=967200 $Y=507100
X963 5430 1 2 5443 DELB $T=969060 426840 1 0 $X=969060 $Y=421420
X964 5441 1 2 5459 DELB $T=973400 527640 0 0 $X=973400 $Y=527260
X965 5436 1 2 5447 DELB $T=975260 406680 1 0 $X=975260 $Y=401260
X966 5377 1 2 5396 DELB $T=975880 487320 0 0 $X=975880 $Y=486940
X967 4909 1 2 4921 DELB $T=978980 487320 1 0 $X=978980 $Y=481900
X968 5471 1 2 5474 DELB $T=980220 507480 1 0 $X=980220 $Y=502060
X969 955 1 2 965 DELB $T=983320 386520 1 0 $X=983320 $Y=381100
X970 5480 1 2 5502 DELB $T=983940 406680 0 0 $X=983940 $Y=406300
X971 5437 1 2 5509 DELB $T=985180 487320 1 0 $X=985180 $Y=481900
X972 5524 1 2 5533 DELB $T=990140 457080 0 0 $X=990140 $Y=456700
X973 5488 1 2 5530 DELB $T=991380 406680 0 0 $X=991380 $Y=406300
X974 5551 1 2 5561 DELB $T=1000680 487320 0 0 $X=1000680 $Y=486940
X975 5523 1 2 5565 DELB $T=1001920 457080 1 0 $X=1001920 $Y=451660
X976 5618 1 2 5626 DELB $T=1008120 416760 0 0 $X=1008120 $Y=416380
X977 5639 1 2 5645 DELB $T=1012460 487320 0 0 $X=1012460 $Y=486940
X978 5660 1 2 5656 DELB $T=1017420 386520 1 0 $X=1017420 $Y=381100
X979 5663 1 2 5617 DELB $T=1018660 497400 1 0 $X=1018660 $Y=491980
X980 5682 1 2 5685 DELB $T=1024240 416760 1 0 $X=1024240 $Y=411340
X981 5686 1 2 5696 DELB $T=1024240 447000 1 0 $X=1024240 $Y=441580
X982 5703 1 2 5705 DELB $T=1028580 436920 0 0 $X=1028580 $Y=436540
X983 5694 1 2 5724 DELB $T=1029200 517560 1 0 $X=1029200 $Y=512140
X984 5719 1 2 5738 DELB $T=1031060 386520 0 0 $X=1031060 $Y=386140
X985 1040 1 2 1048 DELB $T=1032300 497400 1 0 $X=1032300 $Y=491980
X986 5731 1 2 5741 DELB $T=1034780 376440 1 0 $X=1034780 $Y=371020
X987 5702 1 2 5701 DELB $T=1034780 477240 1 0 $X=1034780 $Y=471820
X988 5736 1 2 5756 DELB $T=1034780 507480 0 0 $X=1034780 $Y=507100
X989 5752 1 2 5773 DELB $T=1038500 497400 1 0 $X=1038500 $Y=491980
X990 5707 1 2 5716 DELB $T=1040360 376440 0 0 $X=1040360 $Y=376060
X991 5739 1 2 5757 DELB $T=1041600 396600 1 0 $X=1041600 $Y=391180
X992 5747 1 2 5767 DELB $T=1041600 426840 1 0 $X=1041600 $Y=421420
X993 5774 1 2 5798 DELB $T=1042840 497400 0 0 $X=1042840 $Y=497020
X994 5782 1 2 5806 DELB $T=1045320 426840 0 0 $X=1045320 $Y=426460
X995 5791 1 2 5777 DELB $T=1046560 467160 1 0 $X=1046560 $Y=461740
X996 5797 1 2 5795 DELB $T=1047800 497400 1 0 $X=1047800 $Y=491980
X997 5801 1 2 5794 DELB $T=1048420 396600 1 0 $X=1048420 $Y=391180
X998 5785 1 2 5799 DELB $T=1048420 527640 0 0 $X=1048420 $Y=527260
X999 5820 1 2 5843 DELB $T=1052760 517560 0 0 $X=1052760 $Y=517180
X1000 1070 1 2 5822 DELB $T=1054000 366360 0 0 $X=1054000 $Y=365980
X1001 5826 1 2 5832 DELB $T=1054620 426840 0 0 $X=1054620 $Y=426460
X1002 5841 1 2 5862 DELB $T=1057720 396600 1 0 $X=1057720 $Y=391180
X1003 5813 1 2 5849 DELB $T=1058960 467160 0 0 $X=1058960 $Y=466780
X1004 5869 1 2 5902 DELB $T=1064540 376440 0 0 $X=1064540 $Y=376060
X1005 5870 1 2 5879 DELB $T=1064540 406680 1 0 $X=1064540 $Y=401260
X1006 5885 1 2 5883 DELB $T=1067020 507480 0 0 $X=1067020 $Y=507100
X1007 5850 1 2 5873 DELB $T=1068880 386520 1 0 $X=1068880 $Y=381100
X1008 5835 1 2 5857 DELB $T=1071360 447000 0 0 $X=1071360 $Y=446620
X1009 5928 1 2 5931 DELB $T=1075700 477240 1 0 $X=1075700 $Y=471820
X1010 5937 1 2 5945 DELB $T=1077560 447000 0 0 $X=1077560 $Y=446620
X1011 5909 1 2 5924 DELB $T=1078800 507480 0 0 $X=1078800 $Y=507100
X1012 5955 1 2 5975 DELB $T=1081900 416760 0 0 $X=1081900 $Y=416380
X1013 5956 1 2 5959 DELB $T=1082520 467160 1 0 $X=1082520 $Y=461740
X1014 5958 1 2 5946 DELB $T=1082520 477240 1 0 $X=1082520 $Y=471820
X1015 5960 1 2 5974 DELB $T=1083140 537720 1 0 $X=1083140 $Y=532300
X1016 5890 1 2 5904 DELB $T=1084380 436920 1 0 $X=1084380 $Y=431500
X1017 5979 1 2 6004 DELB $T=1087480 527640 1 0 $X=1087480 $Y=522220
X1018 5986 1 2 6006 DELB $T=1088720 396600 0 0 $X=1088720 $Y=396220
X1019 5997 1 2 6002 DELB $T=1091820 406680 1 0 $X=1091820 $Y=401260
X1020 6008 1 2 6028 DELB $T=1096780 426840 0 0 $X=1096780 $Y=426460
X1021 6046 1 2 6090 DELB $T=1106080 396600 0 0 $X=1106080 $Y=396220
X1022 6054 1 2 6075 DELB $T=1107940 376440 0 0 $X=1107940 $Y=376060
X1023 5983 1 2 6024 DELB $T=1109180 527640 0 0 $X=1109180 $Y=527260
X1024 6038 1 2 6101 DELB $T=1110420 426840 0 0 $X=1110420 $Y=426460
X1025 6076 1 2 6093 DELB $T=1110420 497400 0 0 $X=1110420 $Y=497020
X1026 6095 1 2 6122 DELB $T=1111040 416760 0 0 $X=1111040 $Y=416380
X1027 6013 1 2 6104 DELB $T=1116620 386520 1 0 $X=1116620 $Y=381100
X1028 6056 1 2 6121 DELB $T=1116620 537720 1 0 $X=1116620 $Y=532300
X1029 6078 1 2 6135 DELB $T=1122820 416760 1 0 $X=1122820 $Y=411340
X1030 6109 1 2 6137 DELB $T=1123440 537720 1 0 $X=1123440 $Y=532300
X1031 6069 1 2 6133 DELB $T=1124680 396600 0 0 $X=1124680 $Y=396220
X1032 1721 1 2 1764 DELA $T=311860 376440 0 0 $X=311860 $Y=376060
X1033 1791 1 2 1822 DELA $T=322400 396600 1 0 $X=322400 $Y=391180
X1034 1796 1 2 1820 DELA $T=322400 487320 1 0 $X=322400 $Y=481900
X1035 1803 1 2 1790 DELA $T=323640 426840 0 0 $X=323640 $Y=426460
X1036 1815 1 2 1816 DELA $T=325500 406680 1 0 $X=325500 $Y=401260
X1037 1828 1 2 1812 DELA $T=327980 386520 0 0 $X=327980 $Y=386140
X1038 1845 1 2 1807 DELA $T=330460 406680 1 0 $X=330460 $Y=401260
X1039 117 1 2 1799 DELA $T=331700 436920 0 0 $X=331700 $Y=436540
X1040 1844 1 2 1806 DELA $T=336040 376440 1 0 $X=336040 $Y=371020
X1041 2374 1 2 2410 DELA $T=420980 477240 0 0 $X=420980 $Y=476860
X1042 2375 1 2 2462 DELA $T=429660 497400 0 0 $X=429660 $Y=497020
X1043 2411 1 2 2484 DELA $T=434000 497400 1 0 $X=434000 $Y=491980
X1044 2299 1 2 2390 DELA $T=440820 477240 1 0 $X=440820 $Y=471820
X1045 2212 1 2 2442 DELA $T=445780 477240 1 0 $X=445780 $Y=471820
X1046 2578 1 2 2582 DELA $T=452600 527640 1 0 $X=452600 $Y=522220
X1047 2606 1 2 2618 DELA $T=457560 527640 1 0 $X=457560 $Y=522220
X1048 2621 1 2 2652 DELA $T=461280 416760 0 0 $X=461280 $Y=416380
X1049 2720 1 2 2745 DELA $T=479880 487320 0 0 $X=479880 $Y=486940
X1050 3626 1 2 3656 DELA $T=608840 487320 1 0 $X=608840 $Y=481900
X1051 3641 1 2 3668 DELA $T=610080 527640 1 0 $X=610080 $Y=522220
X1052 3675 1 2 3703 DELA $T=615040 527640 1 0 $X=615040 $Y=522220
X1053 3765 1 2 3797 DELA $T=631160 467160 1 0 $X=631160 $Y=461740
X1054 3804 1 2 3824 DELA $T=636740 447000 0 0 $X=636740 $Y=446620
X1055 3841 1 2 3869 DELA $T=643560 497400 0 0 $X=643560 $Y=497020
X1056 3928 1 2 3960 DELA $T=657820 426840 0 0 $X=657820 $Y=426460
X1057 3952 1 2 3979 DELA $T=662160 426840 1 0 $X=662160 $Y=421420
X1058 3990 1 2 4017 DELA $T=670220 426840 0 0 $X=670220 $Y=426460
X1059 3999 1 2 4029 DELA $T=672080 436920 1 0 $X=672080 $Y=431500
X1060 4021 1 2 4044 DELA $T=675180 426840 0 0 $X=675180 $Y=426460
X1061 4039 1 2 4063 DELA $T=678280 497400 0 0 $X=678280 $Y=497020
X1062 4060 1 2 4075 DELA $T=681380 386520 0 0 $X=681380 $Y=386140
X1063 4064 1 2 4085 DELA $T=683240 497400 0 0 $X=683240 $Y=497020
X1064 4079 1 2 4102 DELA $T=686340 386520 0 0 $X=686340 $Y=386140
X1065 547 1 2 553 DELA $T=686960 537720 1 0 $X=686960 $Y=532300
X1066 4095 1 2 4117 DELA $T=690060 426840 0 0 $X=690060 $Y=426460
X1067 4107 1 2 4125 DELA $T=691300 386520 0 0 $X=691300 $Y=386140
X1068 4129 1 2 4130 DELA $T=696260 386520 0 0 $X=696260 $Y=386140
X1069 4287 1 2 4283 DELA $T=728500 416760 0 0 $X=728500 $Y=416380
X1070 4294 1 2 4327 DELA $T=730980 376440 0 0 $X=730980 $Y=376060
X1071 4758 1 2 4767 DELA $T=831420 457080 1 0 $X=831420 $Y=451660
X1072 5108 1 2 5136 DELA $T=901480 447000 0 0 $X=901480 $Y=446620
X1073 5128 1 2 5168 DELA $T=906440 447000 0 0 $X=906440 $Y=446620
X1074 5139 1 2 5172 DELA $T=907060 507480 0 0 $X=907060 $Y=507100
X1075 5260 1 2 5253 DELA $T=936820 447000 1 0 $X=936820 $Y=441580
X1076 5302 1 2 5313 DELA $T=942400 376440 1 0 $X=942400 $Y=371020
X1077 882 1 2 894 DELA $T=944260 537720 1 0 $X=944260 $Y=532300
X1078 5267 1 2 5210 DELA $T=946120 457080 0 0 $X=946120 $Y=456700
X1079 5234 1 2 5157 DELA $T=952940 426840 0 0 $X=952940 $Y=426460
X1080 914 1 2 921 DELA $T=957280 527640 0 0 $X=957280 $Y=527260
X1081 919 1 2 925 DELA $T=961000 396600 1 0 $X=961000 $Y=391180
X1082 5123 1 2 5150 DELA $T=966580 426840 0 0 $X=966580 $Y=426460
X1083 5389 1 2 5406 DELA $T=969060 477240 0 0 $X=969060 $Y=476860
X1084 928 1 2 934 DELA $T=971540 386520 0 0 $X=971540 $Y=386140
X1085 5280 1 2 5350 DELA $T=972160 497400 1 0 $X=972160 $Y=491980
X1086 5448 1 2 5465 DELA $T=983320 396600 1 0 $X=983320 $Y=391180
X1087 5496 1 2 5521 DELA $T=988280 386520 1 0 $X=988280 $Y=381100
X1088 5446 1 2 5494 DELA $T=990760 497400 0 0 $X=990760 $Y=497020
X1089 5525 1 2 5522 DELA $T=994480 447000 1 0 $X=994480 $Y=441580
X1090 5528 1 2 5534 DELA $T=995720 497400 0 0 $X=995720 $Y=497020
X1091 5564 1 2 5600 DELA $T=999440 447000 1 0 $X=999440 $Y=441580
X1092 5552 1 2 5576 DELA $T=1000680 497400 0 0 $X=1000680 $Y=497020
X1093 5541 1 2 5569 DELA $T=1019900 467160 1 0 $X=1019900 $Y=461740
X1094 5706 1 2 5746 DELA $T=1032920 527640 1 0 $X=1032920 $Y=522220
X1095 5844 1 2 5819 DELA $T=1063920 467160 0 0 $X=1063920 $Y=466780
X1096 1223 23 30 2 1 1205 QDFFRBN $T=225060 527640 0 0 $X=225060 $Y=527260
X1097 1256 23 30 2 1 1234 QDFFRBN $T=230020 537720 1 0 $X=230020 $Y=532300
X1098 40 23 30 2 1 47 QDFFRBN $T=243660 537720 1 0 $X=243660 $Y=532300
X1099 1735 23 1787 2 1 108 QDFFRBN $T=313100 457080 0 0 $X=313100 $Y=456700
X1100 1754 23 1787 2 1 1796 QDFFRBN $T=314960 477240 1 0 $X=314960 $Y=471820
X1101 1762 23 1805 2 1 117 QDFFRBN $T=315580 436920 1 0 $X=315580 $Y=431500
X1102 1779 114 118 2 1 1844 QDFFRBN $T=319300 366360 0 0 $X=319300 $Y=365980
X1103 1782 23 1787 2 1 107 QDFFRBN $T=319300 447000 0 0 $X=319300 $Y=446620
X1104 1792 114 118 2 1 1828 QDFFRBN $T=321780 386520 1 0 $X=321780 $Y=381100
X1105 1793 23 1805 2 1 1840 QDFFRBN $T=321780 416760 0 0 $X=321780 $Y=416380
X1106 1809 114 1805 2 1 1803 QDFFRBN $T=323640 416760 1 0 $X=323640 $Y=411340
X1107 1810 114 1853 2 1 1721 QDFFRBN $T=324260 376440 1 0 $X=324260 $Y=371020
X1108 1813 114 1805 2 1 1845 QDFFRBN $T=326740 396600 0 0 $X=326740 $Y=396220
X1109 1827 114 1805 2 1 1815 QDFFRBN $T=326740 406680 0 0 $X=326740 $Y=406300
X1110 1842 23 1787 2 1 125 QDFFRBN $T=329840 487320 1 0 $X=329840 $Y=481900
X1111 1846 23 1787 2 1 1862 QDFFRBN $T=330460 497400 1 0 $X=330460 $Y=491980
X1112 1859 114 1853 2 1 1791 QDFFRBN $T=332940 396600 1 0 $X=332940 $Y=391180
X1113 2394 231 1853 2 1 2299 QDFFRBN $T=434620 447000 1 180 $X=422840 $Y=446620
X1114 2436 231 2433 2 1 2374 QDFFRBN $T=437720 477240 1 180 $X=425940 $Y=476860
X1115 2439 231 2433 2 1 2402 QDFFRBN $T=438960 457080 0 180 $X=427180 $Y=451660
X1116 2441 231 2433 2 1 2212 QDFFRBN $T=441440 457080 1 180 $X=429660 $Y=456700
X1117 2494 231 2433 2 1 2399 QDFFRBN $T=442680 467160 0 180 $X=430900 $Y=461740
X1118 2483 231 2488 2 1 2411 QDFFRBN $T=447020 487320 0 180 $X=435240 $Y=481900
X1119 2506 231 2488 2 1 2375 QDFFRBN $T=450740 497400 0 180 $X=438960 $Y=491980
X1120 250 253 256 2 1 246 QDFFRBN $T=443300 537720 1 0 $X=443300 $Y=532300
X1121 2538 231 2583 2 1 2516 QDFFRBN $T=445780 507480 1 0 $X=445780 $Y=502060
X1122 2553 231 256 2 1 2372 QDFFRBN $T=447640 517560 1 0 $X=447640 $Y=512140
X1123 2582 231 2583 2 1 2613 QDFFRBN $T=453220 497400 0 0 $X=453220 $Y=497020
X1124 2596 231 2570 2 1 2666 QDFFRBN $T=456320 477240 1 0 $X=456320 $Y=471820
X1125 2663 231 2583 2 1 2675 QDFFRBN $T=466860 497400 0 0 $X=466860 $Y=497020
X1126 2654 231 2583 2 1 2606 QDFFRBN $T=469340 507480 1 0 $X=469340 $Y=502060
X1127 2745 231 2570 2 1 2611 QDFFRBN $T=481740 477240 0 180 $X=469960 $Y=471820
X1128 2692 231 2735 2 1 2763 QDFFRBN $T=471200 416760 0 0 $X=471200 $Y=416380
X1129 2694 231 2646 2 1 2788 QDFFRBN $T=471820 426840 1 0 $X=471820 $Y=421420
X1130 2718 231 2646 2 1 2789 QDFFRBN $T=475540 436920 1 0 $X=475540 $Y=431500
X1131 2728 231 2570 2 1 2806 QDFFRBN $T=477400 467160 0 0 $X=477400 $Y=466780
X1132 2732 231 2735 2 1 2800 QDFFRBN $T=478640 396600 0 0 $X=478640 $Y=396220
X1133 2740 231 2646 2 1 2784 QDFFRBN $T=479260 447000 0 0 $X=479260 $Y=446620
X1134 2744 231 2735 2 1 2816 QDFFRBN $T=479880 406680 0 0 $X=479880 $Y=406300
X1135 2755 231 2735 2 1 2815 QDFFRBN $T=481120 406680 1 0 $X=481120 $Y=401260
X1136 2762 231 2735 2 1 2821 QDFFRBN $T=482980 396600 1 0 $X=482980 $Y=391180
X1137 2765 231 2646 2 1 2824 QDFFRBN $T=482980 447000 1 0 $X=482980 $Y=441580
X1138 2766 231 2570 2 1 2726 QDFFRBN $T=482980 467160 1 0 $X=482980 $Y=461740
X1139 2767 231 2570 2 1 2835 QDFFRBN $T=483600 477240 1 0 $X=483600 $Y=471820
X1140 2768 231 2749 2 1 2796 QDFFRBN $T=483600 507480 1 0 $X=483600 $Y=502060
X1141 2798 231 2813 2 1 2874 QDFFRBN $T=489180 386520 1 0 $X=489180 $Y=381100
X1142 2807 231 2749 2 1 2858 QDFFRBN $T=490420 507480 0 0 $X=490420 $Y=507100
X1143 2829 231 320 2 1 334 QDFFRBN $T=494760 366360 0 0 $X=494760 $Y=365980
X1144 2927 231 2813 2 1 2833 QDFFRBN $T=507160 396600 0 180 $X=495380 $Y=391180
X1145 2868 231 2749 2 1 324 QDFFRBN $T=507160 527640 0 180 $X=495380 $Y=522220
X1146 2840 231 320 2 1 332 QDFFRBN $T=496000 376440 1 0 $X=496000 $Y=371020
X1147 2841 231 320 2 1 2883 QDFFRBN $T=496000 376440 0 0 $X=496000 $Y=376060
X1148 2913 231 2813 2 1 2843 QDFFRBN $T=508400 386520 1 180 $X=496620 $Y=386140
X1149 2873 231 2825 2 1 2864 QDFFRBN $T=510880 457080 1 180 $X=499100 $Y=456700
X1150 3021 231 320 2 1 331 QDFFRBN $T=520180 366360 1 180 $X=508400 $Y=365980
X1151 3062 231 2783 2 1 2974 QDFFRBN $T=525760 426840 0 180 $X=513980 $Y=421420
X1152 3156 231 2783 2 1 3074 QDFFRBN $T=536920 426840 1 180 $X=525140 $Y=426460
X1153 3057 231 2749 2 1 349 QDFFRBN $T=525760 527640 0 0 $X=525760 $Y=527260
X1154 3090 231 2749 2 1 351 QDFFRBN $T=525760 537720 1 0 $X=525760 $Y=532300
X1155 3171 231 2783 2 1 3094 QDFFRBN $T=538780 426840 0 180 $X=527000 $Y=421420
X1156 3199 231 2825 2 1 3126 QDFFRBN $T=541880 467160 1 180 $X=530100 $Y=466780
X1157 3160 231 2825 2 1 2830 QDFFRBN $T=534440 467160 1 0 $X=534440 $Y=461740
X1158 3210 231 2783 2 1 3163 QDFFRBN $T=549940 426840 1 180 $X=538160 $Y=426460
X1159 3192 231 3240 2 1 3054 QDFFRBN $T=539400 527640 0 0 $X=539400 $Y=527260
X1160 3265 231 2783 2 1 3153 QDFFRBN $T=551800 426840 0 180 $X=540020 $Y=421420
X1161 3164 231 2825 2 1 3287 QDFFRBN $T=541260 477240 1 0 $X=541260 $Y=471820
X1162 3129 231 3240 2 1 406 QDFFRBN $T=547460 517560 0 0 $X=547460 $Y=517180
X1163 3260 231 3288 2 1 3323 QDFFRBN $T=556760 527640 0 0 $X=556760 $Y=527260
X1164 3333 231 3288 2 1 3394 QDFFRBN $T=561100 517560 0 0 $X=561100 $Y=517180
X1165 3918 3926 3948 2 1 3961 QDFFRBN $T=654720 487320 0 0 $X=654720 $Y=486940
X1166 3935 518 3981 2 1 3983 QDFFRBN $T=658440 507480 0 0 $X=658440 $Y=507100
X1167 3943 3926 3986 2 1 4015 QDFFRBN $T=659680 457080 0 0 $X=659680 $Y=456700
X1168 3944 3926 3986 2 1 3993 QDFFRBN $T=659680 467160 1 0 $X=659680 $Y=461740
X1169 3945 518 513 2 1 529 QDFFRBN $T=659680 537720 1 0 $X=659680 $Y=532300
X1170 3989 3926 3948 2 1 3947 QDFFRBN $T=672080 487320 0 180 $X=660300 $Y=481900
X1171 3958 518 3948 2 1 3927 QDFFRBN $T=661540 507480 1 0 $X=661540 $Y=502060
X1172 3964 3926 3986 2 1 3980 QDFFRBN $T=662160 447000 0 0 $X=662160 $Y=446620
X1173 3965 3926 3986 2 1 3626 QDFFRBN $T=662160 477240 0 0 $X=662160 $Y=476860
X1174 3998 518 3972 2 1 4046 QDFFRBN $T=671460 517560 0 0 $X=671460 $Y=517180
X1175 4006 518 3972 2 1 3675 QDFFRBN $T=672700 507480 0 0 $X=672700 $Y=507100
X1176 4023 518 3948 2 1 3801 QDFFRBN $T=675180 507480 1 0 $X=675180 $Y=502060
X1177 4011 518 3972 2 1 3707 QDFFRBN $T=675800 527640 1 0 $X=675800 $Y=522220
X1178 4028 541 4056 2 1 4052 QDFFRBN $T=676420 426840 1 0 $X=676420 $Y=421420
X1179 4030 3926 4069 2 1 3954 QDFFRBN $T=676420 447000 0 0 $X=676420 $Y=446620
X1180 4031 3926 3981 2 1 4013 QDFFRBN $T=676420 487320 1 0 $X=676420 $Y=481900
X1181 4035 3926 4056 2 1 3928 QDFFRBN $T=677040 436920 1 0 $X=677040 $Y=431500
X1182 4084 3926 3948 2 1 4004 QDFFRBN $T=689440 487320 1 180 $X=677660 $Y=486940
X1183 4040 3926 4056 2 1 4104 QDFFRBN $T=678280 436920 0 0 $X=678280 $Y=436540
X1184 4042 3926 4033 2 1 4096 QDFFRBN $T=678900 467160 0 0 $X=678900 $Y=466780
X1185 550 518 544 2 1 4054 QDFFRBN $T=691920 527640 1 180 $X=680140 $Y=527260
X1186 4065 3926 4033 2 1 4062 QDFFRBN $T=683240 467160 1 0 $X=683240 $Y=461740
X1187 4067 541 4111 2 1 4107 QDFFRBN $T=683860 396600 0 0 $X=683860 $Y=396220
X1188 4078 541 4056 2 1 4133 QDFFRBN $T=685720 416760 1 0 $X=685720 $Y=411340
X1189 4082 541 4111 2 1 4129 QDFFRBN $T=686960 406680 0 0 $X=686960 $Y=406300
X1190 4083 3926 4033 2 1 3999 QDFFRBN $T=686960 457080 1 0 $X=686960 $Y=451660
X1191 4086 518 4033 2 1 4039 QDFFRBN $T=688200 507480 1 0 $X=688200 $Y=502060
X1192 4094 541 4136 2 1 4079 QDFFRBN $T=689440 396600 1 0 $X=689440 $Y=391180
X1193 4145 518 4080 2 1 4098 QDFFRBN $T=701840 517560 0 180 $X=690060 $Y=512140
X1194 4108 541 4136 2 1 4060 QDFFRBN $T=691300 386520 1 0 $X=691300 $Y=381100
X1195 4162 3926 4033 2 1 4064 QDFFRBN $T=703080 487320 1 180 $X=691300 $Y=486940
X1196 4110 518 4080 2 1 4109 QDFFRBN $T=691300 527640 1 0 $X=691300 $Y=522220
X1197 4193 3926 4156 2 1 4137 QDFFRBN $T=709280 467160 0 180 $X=697500 $Y=461740
X1198 4147 3926 4069 2 1 4160 QDFFRBN $T=698120 447000 1 0 $X=698120 $Y=441580
X1199 4189 3926 3981 2 1 4144 QDFFRBN $T=709900 487320 0 180 $X=698120 $Y=481900
X1200 4157 3926 4156 2 1 4150 QDFFRBN $T=699980 457080 0 0 $X=699980 $Y=456700
X1201 4158 541 572 2 1 4143 QDFFRBN $T=700600 376440 1 0 $X=700600 $Y=371020
X1202 4164 541 4111 2 1 4020 QDFFRBN $T=701840 406680 0 0 $X=701840 $Y=406300
X1203 4169 541 572 2 1 4113 QDFFRBN $T=702460 366360 0 0 $X=702460 $Y=365980
X1204 4175 3926 4156 2 1 3841 QDFFRBN $T=704940 487320 0 0 $X=704940 $Y=486940
X1205 4241 3926 4069 2 1 4177 QDFFRBN $T=717340 426840 1 180 $X=705560 $Y=426460
X1206 4186 541 4111 2 1 4176 QDFFRBN $T=706180 406680 1 0 $X=706180 $Y=401260
X1207 4183 541 4111 2 1 4191 QDFFRBN $T=706800 396600 0 0 $X=706800 $Y=396220
X1208 4190 518 4080 2 1 584 QDFFRBN $T=706800 527640 1 0 $X=706800 $Y=522220
X1209 4180 518 4080 2 1 3811 QDFFRBN $T=707420 517560 0 0 $X=707420 $Y=517180
X1210 4232 3926 4069 2 1 4072 QDFFRBN $T=719820 436920 0 180 $X=708040 $Y=431500
X1211 4233 3926 4156 2 1 3952 QDFFRBN $T=719820 457080 0 180 $X=708040 $Y=451660
X1212 4198 518 4226 2 1 4209 QDFFRBN $T=708660 507480 1 0 $X=708660 $Y=502060
X1213 4185 518 4080 2 1 3695 QDFFRBN $T=722300 517560 0 180 $X=710520 $Y=512140
X1214 4201 3926 4237 2 1 4212 QDFFRBN $T=711140 487320 1 0 $X=711140 $Y=481900
X1215 4207 3926 4156 2 1 3765 QDFFRBN $T=723540 467160 0 180 $X=711760 $Y=461740
X1216 4278 541 572 2 1 4221 QDFFRBN $T=727880 386520 0 180 $X=716100 $Y=381100
X1217 4257 541 4223 2 1 4222 QDFFRBN $T=727880 406680 1 180 $X=716100 $Y=406300
X1218 4266 541 572 2 1 4224 QDFFRBN $T=728500 366360 1 180 $X=716720 $Y=365980
X1219 4273 541 572 2 1 4227 QDFFRBN $T=729120 396600 0 180 $X=717340 $Y=391180
X1220 4234 518 4226 2 1 587 QDFFRBN $T=717960 537720 1 0 $X=717960 $Y=532300
X1221 4236 3926 4237 2 1 4217 QDFFRBN $T=718580 487320 0 0 $X=718580 $Y=486940
X1222 4275 518 4252 2 1 4235 QDFFRBN $T=730360 497400 1 180 $X=718580 $Y=497020
X1223 4244 518 4226 2 1 4300 QDFFRBN $T=720440 527640 1 0 $X=720440 $Y=522220
X1224 4250 3926 4223 2 1 4287 QDFFRBN $T=721060 426840 1 0 $X=721060 $Y=421420
X1225 4318 3926 4237 2 1 4260 QDFFRBN $T=735320 467160 0 180 $X=723540 $Y=461740
X1226 4261 3926 4237 2 1 4247 QDFFRBN $T=723540 477240 0 0 $X=723540 $Y=476860
X1227 4267 518 4226 2 1 4296 QDFFRBN $T=724160 517560 1 0 $X=724160 $Y=512140
X1228 4277 541 596 2 1 603 QDFFRBN $T=725400 376440 1 0 $X=725400 $Y=371020
X1229 4330 3926 4223 2 1 4021 QDFFRBN $T=737800 416760 0 180 $X=726020 $Y=411340
X1230 4279 3926 4303 2 1 4312 QDFFRBN $T=726020 447000 0 0 $X=726020 $Y=446620
X1231 4286 541 4323 2 1 600 QDFFRBN $T=727260 396600 0 0 $X=727260 $Y=396220
X1232 4350 541 596 2 1 4302 QDFFRBN $T=743380 366360 1 180 $X=731600 $Y=365980
X1233 4347 541 4323 2 1 4294 QDFFRBN $T=743380 396600 0 180 $X=731600 $Y=391180
X1234 4311 518 4226 2 1 3742 QDFFRBN $T=732220 517560 0 0 $X=732220 $Y=517180
X1235 4362 612 4252 2 1 4325 QDFFRBN $T=746480 497400 0 180 $X=734700 $Y=491980
X1236 4361 3926 4237 2 1 4280 QDFFRBN $T=747100 467160 0 180 $X=735320 $Y=461740
X1237 4345 3926 4338 2 1 4326 QDFFRBN $T=747100 477240 1 180 $X=735320 $Y=476860
X1238 4366 612 4226 2 1 4329 QDFFRBN $T=747100 507480 1 180 $X=735320 $Y=507100
X1239 4333 3926 4323 2 1 621 QDFFRBN $T=736560 406680 0 0 $X=736560 $Y=406300
X1240 4349 3926 4338 2 1 4309 QDFFRBN $T=748960 487320 0 180 $X=737180 $Y=481900
X1241 4334 518 614 2 1 4293 QDFFRBN $T=737180 527640 0 0 $X=737180 $Y=527260
X1242 4378 3926 4223 2 1 601 QDFFRBN $T=749580 416760 0 180 $X=737800 $Y=411340
X1243 4337 3926 4303 2 1 4352 QDFFRBN $T=737800 436920 0 0 $X=737800 $Y=436540
X1244 4342 3926 4377 2 1 4364 QDFFRBN $T=739660 426840 0 0 $X=739660 $Y=426460
X1245 4346 541 4323 2 1 4373 QDFFRBN $T=740280 386520 0 0 $X=740280 $Y=386140
X1246 4355 518 614 2 1 4270 QDFFRBN $T=742760 527640 1 0 $X=742760 $Y=522220
X1247 4417 628 596 2 1 4367 QDFFRBN $T=757640 376440 0 180 $X=745860 $Y=371020
X1248 4360 541 4408 2 1 4374 QDFFRBN $T=746480 396600 1 0 $X=746480 $Y=391180
X1249 4421 628 4323 2 1 4369 QDFFRBN $T=758260 406680 0 180 $X=746480 $Y=401260
X1250 4375 612 4252 2 1 3893 QDFFRBN $T=747100 517560 1 0 $X=747100 $Y=512140
X1251 4379 612 4338 2 1 4420 QDFFRBN $T=747720 497400 0 0 $X=747720 $Y=497020
X1252 4386 612 4252 2 1 3739 QDFFRBN $T=748960 507480 1 0 $X=748960 $Y=502060
X1253 4413 3926 4404 2 1 4395 QDFFRBN $T=763220 457080 1 180 $X=751440 $Y=456700
X1254 4397 3926 4338 2 1 3874 QDFFRBN $T=751440 477240 0 0 $X=751440 $Y=476860
X1255 4445 3926 4404 2 1 3970 QDFFRBN $T=763840 467160 0 180 $X=752060 $Y=461740
X1256 4451 628 4408 2 1 4403 QDFFRBN $T=764460 386520 0 180 $X=752680 $Y=381100
X1257 4435 3926 4338 2 1 3667 QDFFRBN $T=766320 477240 0 180 $X=754540 $Y=471820
X1258 4432 612 614 2 1 3641 QDFFRBN $T=768800 527640 1 180 $X=757020 $Y=527260
X1259 4454 3926 4431 2 1 3985 QDFFRBN $T=769420 436920 1 180 $X=757640 $Y=436540
X1260 4425 3926 4404 2 1 4480 QDFFRBN $T=757640 447000 0 0 $X=757640 $Y=446620
X1261 4427 628 4465 2 1 4484 QDFFRBN $T=758260 376440 1 0 $X=758260 $Y=371020
X1262 4428 3926 4377 2 1 4471 QDFFRBN $T=758260 436920 1 0 $X=758260 $Y=431500
X1263 643 612 614 2 1 635 QDFFRBN $T=771280 537720 0 180 $X=759500 $Y=532300
X1264 4434 3926 4377 2 1 4422 QDFFRBN $T=760120 416760 0 0 $X=760120 $Y=416380
X1265 4458 3926 4494 2 1 4473 QDFFRBN $T=763840 497400 1 0 $X=763840 $Y=491980
X1266 4468 628 4465 2 1 4499 QDFFRBN $T=765700 406680 1 0 $X=765700 $Y=401260
X1267 4469 612 4483 2 1 648 QDFFRBN $T=765700 527640 1 0 $X=765700 $Y=522220
X1268 4455 3926 4481 2 1 4447 QDFFRBN $T=766320 467160 1 0 $X=766320 $Y=461740
X1269 4493 3926 4481 2 1 4460 QDFFRBN $T=778720 477240 1 180 $X=766940 $Y=476860
X1270 4532 628 4408 2 1 4476 QDFFRBN $T=779960 386520 1 180 $X=768180 $Y=386140
X1271 4488 3926 4431 2 1 4314 QDFFRBN $T=770040 426840 0 0 $X=770040 $Y=426460
X1272 4522 3926 4481 2 1 3919 QDFFRBN $T=782440 457080 1 180 $X=770660 $Y=456700
X1273 4542 628 4465 2 1 4490 QDFFRBN $T=783060 376440 0 180 $X=771280 $Y=371020
X1274 4500 3926 4539 2 1 4440 QDFFRBN $T=771900 457080 1 0 $X=771900 $Y=451660
X1275 4549 628 4431 2 1 4502 QDFFRBN $T=784300 436920 0 180 $X=772520 $Y=431500
X1276 657 612 614 2 1 646 QDFFRBN $T=785540 537720 0 180 $X=773760 $Y=532300
X1277 4561 628 4408 2 1 4519 QDFFRBN $T=788020 396600 0 180 $X=776240 $Y=391180
X1278 650 628 658 2 1 660 QDFFRBN $T=777480 366360 0 0 $X=777480 $Y=365980
X1279 4536 3926 4539 2 1 4571 QDFFRBN $T=778720 477240 1 0 $X=778720 $Y=471820
X1280 4495 612 659 2 1 3551 QDFFRBN $T=778720 527640 1 0 $X=778720 $Y=522220
X1281 4547 628 4465 2 1 4489 QDFFRBN $T=791120 406680 0 180 $X=779340 $Y=401260
X1282 4557 3926 4539 2 1 4533 QDFFRBN $T=792360 467160 0 180 $X=780580 $Y=461740
X1283 4504 3926 4539 2 1 3857 QDFFRBN $T=780580 477240 0 0 $X=780580 $Y=476860
X1284 4531 612 659 2 1 3587 QDFFRBN $T=780580 517560 1 0 $X=780580 $Y=512140
X1285 4543 628 4570 2 1 4568 QDFFRBN $T=781200 416760 1 0 $X=781200 $Y=411340
X1286 4517 612 4494 2 1 4479 QDFFRBN $T=781820 507480 0 0 $X=781820 $Y=507100
X1287 4552 612 4494 2 1 4419 QDFFRBN $T=782440 497400 0 0 $X=782440 $Y=497020
X1288 4576 628 4465 2 1 4527 QDFFRBN $T=794840 376440 0 180 $X=783060 $Y=371020
X1289 4559 628 4431 2 1 4535 QDFFRBN $T=794840 426840 1 180 $X=783060 $Y=426460
X1290 4553 3926 4481 2 1 4579 QDFFRBN $T=783060 457080 0 0 $X=783060 $Y=456700
X1291 4558 4560 4481 2 1 4556 QDFFRBN $T=783680 447000 1 0 $X=783680 $Y=441580
X1292 4526 4560 4494 2 1 3784 QDFFRBN $T=796700 487320 1 180 $X=784920 $Y=486940
X1293 4563 628 4591 2 1 4583 QDFFRBN $T=786780 396600 0 0 $X=786780 $Y=396220
X1294 4565 628 4591 2 1 4601 QDFFRBN $T=787400 386520 0 0 $X=787400 $Y=386140
X1295 4587 612 659 2 1 4567 QDFFRBN $T=800420 537720 0 180 $X=788640 $Y=532300
X1296 4618 628 658 2 1 4569 QDFFRBN $T=801040 366360 1 180 $X=789260 $Y=365980
X1297 4585 4560 4626 2 1 4645 QDFFRBN $T=792980 487320 1 0 $X=792980 $Y=481900
X1298 4615 612 659 2 1 4548 QDFFRBN $T=804760 517560 1 180 $X=792980 $Y=517180
X1299 4594 4560 4626 2 1 4640 QDFFRBN $T=794840 457080 0 0 $X=794840 $Y=456700
X1300 4595 4560 4539 2 1 4620 QDFFRBN $T=794840 477240 0 0 $X=794840 $Y=476860
X1301 4600 612 4642 2 1 4643 QDFFRBN $T=795460 517560 1 0 $X=795460 $Y=512140
X1302 4624 628 4570 2 1 4592 QDFFRBN $T=808480 426840 1 180 $X=796700 $Y=426460
X1303 4619 628 4570 2 1 667 QDFFRBN $T=809100 426840 0 180 $X=797320 $Y=421420
X1304 4669 4560 4494 2 1 4612 QDFFRBN $T=809720 497400 0 180 $X=797940 $Y=491980
X1305 4609 4560 4626 2 1 4580 QDFFRBN $T=798560 447000 1 0 $X=798560 $Y=441580
X1306 4613 612 4642 2 1 4681 QDFFRBN $T=799800 527640 1 0 $X=799800 $Y=522220
X1307 4627 628 4670 2 1 669 QDFFRBN $T=801040 386520 0 0 $X=801040 $Y=386140
X1308 4647 612 4642 2 1 685 QDFFRBN $T=804140 537720 1 0 $X=804140 $Y=532300
X1309 4629 628 4570 2 1 675 QDFFRBN $T=816540 416760 1 180 $X=804760 $Y=416380
X1310 4686 628 4670 2 1 4602 QDFFRBN $T=817160 366360 1 180 $X=805380 $Y=365980
X1311 4675 628 4591 2 1 4646 QDFFRBN $T=818400 396600 1 180 $X=806620 $Y=396220
X1312 4696 628 4591 2 1 4637 QDFFRBN $T=819640 416760 0 180 $X=807860 $Y=411340
X1313 4711 628 4670 2 1 668 QDFFRBN $T=821500 396600 0 180 $X=809720 $Y=391180
X1314 4680 628 4670 2 1 4691 QDFFRBN $T=810340 386520 1 0 $X=810340 $Y=381100
X1315 4699 628 591 2 1 4672 QDFFRBN $T=822120 426840 1 180 $X=810340 $Y=426460
X1316 4689 4560 4642 2 1 3844 QDFFRBN $T=822120 517560 0 180 $X=810340 $Y=512140
X1317 4692 4560 4704 2 1 676 QDFFRBN $T=824600 447000 0 180 $X=812820 $Y=441580
X1318 4687 4560 4626 2 1 681 QDFFRBN $T=825220 457080 0 180 $X=813440 $Y=451660
X1319 4665 4560 4719 2 1 677 QDFFRBN $T=813440 497400 1 0 $X=813440 $Y=491980
X1320 4677 4560 4704 2 1 4659 QDFFRBN $T=825840 436920 1 180 $X=814060 $Y=436540
X1321 4688 4560 4626 2 1 4656 QDFFRBN $T=825840 467160 0 180 $X=814060 $Y=461740
X1322 4700 4560 4722 2 1 4733 QDFFRBN $T=814680 477240 1 0 $X=814680 $Y=471820
X1323 4684 4560 4626 2 1 4673 QDFFRBN $T=826460 477240 1 180 $X=814680 $Y=476860
X1324 4703 628 4670 2 1 4735 QDFFRBN $T=815300 376440 1 0 $X=815300 $Y=371020
X1325 4706 4560 4722 2 1 4663 QDFFRBN $T=815920 467160 0 0 $X=815920 $Y=466780
X1326 4715 4560 4719 2 1 4653 QDFFRBN $T=818400 507480 1 0 $X=818400 $Y=502060
X1327 691 696 698 2 1 703 QDFFRBN $T=818400 537720 1 0 $X=818400 $Y=532300
X1328 4716 628 4717 2 1 673 QDFFRBN $T=819020 416760 0 0 $X=819020 $Y=416380
X1329 4709 4560 4722 2 1 4690 QDFFRBN $T=830800 487320 1 180 $X=819020 $Y=486940
X1330 4713 4560 4719 2 1 4698 QDFFRBN $T=831420 497400 1 180 $X=819640 $Y=497020
X1331 4714 696 4642 2 1 4694 QDFFRBN $T=831420 527640 1 180 $X=819640 $Y=527260
X1332 4718 628 4743 2 1 4772 QDFFRBN $T=820260 396600 0 0 $X=820260 $Y=396220
X1333 4723 628 4717 2 1 4750 QDFFRBN $T=822120 406680 0 0 $X=822120 $Y=406300
X1334 4724 628 4717 2 1 706 QDFFRBN $T=822120 426840 1 0 $X=822120 $Y=421420
X1335 4727 628 4756 2 1 4770 QDFFRBN $T=823360 386520 0 0 $X=823360 $Y=386140
X1336 4720 4560 4719 2 1 4012 QDFFRBN $T=835140 527640 0 180 $X=823360 $Y=522220
X1337 4760 4560 4719 2 1 4729 QDFFRBN $T=835760 507480 1 180 $X=823980 $Y=507100
X1338 4740 4560 4751 2 1 4758 QDFFRBN $T=826460 457080 0 0 $X=826460 $Y=456700
X1339 4792 4560 4722 2 1 4738 QDFFRBN $T=838240 497400 0 180 $X=826460 $Y=491980
X1340 4745 4560 4787 2 1 726 QDFFRBN $T=828320 517560 0 0 $X=828320 $Y=517180
X1341 4748 4560 4742 2 1 4766 QDFFRBN $T=828940 436920 0 0 $X=828940 $Y=436540
X1342 4826 4560 4722 2 1 4763 QDFFRBN $T=845060 467160 1 180 $X=833280 $Y=466780
X1343 4802 696 698 2 1 4769 QDFFRBN $T=845680 527640 1 180 $X=833900 $Y=527260
X1344 4788 718 4743 2 1 4784 QDFFRBN $T=836380 406680 0 0 $X=836380 $Y=406300
X1345 4786 718 4743 2 1 714 QDFFRBN $T=848160 426840 0 180 $X=836380 $Y=421420
X1346 4789 4560 4751 2 1 739 QDFFRBN $T=836380 457080 1 0 $X=836380 $Y=451660
X1347 4798 4560 4787 2 1 4835 QDFFRBN $T=838240 507480 0 0 $X=838240 $Y=507100
X1348 4803 718 4742 2 1 4816 QDFFRBN $T=838860 436920 1 0 $X=838860 $Y=431500
X1349 4840 4560 4751 2 1 4800 QDFFRBN $T=850640 457080 1 180 $X=838860 $Y=456700
X1350 4804 4560 4768 2 1 4801 QDFFRBN $T=838860 477240 0 0 $X=838860 $Y=476860
X1351 4807 4560 4787 2 1 4744 QDFFRBN $T=840100 497400 1 0 $X=840100 $Y=491980
X1352 4850 718 4743 2 1 4808 QDFFRBN $T=852500 396600 1 180 $X=840720 $Y=396220
X1353 4810 4560 4787 2 1 748 QDFFRBN $T=841340 517560 0 0 $X=841340 $Y=517180
X1354 4813 718 4756 2 1 749 QDFFRBN $T=841960 376440 0 0 $X=841960 $Y=376060
X1355 4888 4560 4742 2 1 4836 QDFFRBN $T=859320 436920 1 180 $X=847540 $Y=436540
X1356 4837 4560 4787 2 1 4889 QDFFRBN $T=847540 517560 1 0 $X=847540 $Y=512140
X1357 4890 696 4787 2 1 740 QDFFRBN $T=859320 527640 0 180 $X=847540 $Y=522220
X1358 4842 718 4756 2 1 4881 QDFFRBN $T=849400 386520 0 0 $X=849400 $Y=386140
X1359 4904 718 4845 2 1 4843 QDFFRBN $T=861800 426840 0 180 $X=850020 $Y=421420
X1360 4847 4560 4863 2 1 4817 QDFFRBN $T=850020 447000 1 0 $X=850020 $Y=441580
X1361 4848 4560 4863 2 1 4909 QDFFRBN $T=850020 457080 1 0 $X=850020 $Y=451660
X1362 4851 718 4893 2 1 4900 QDFFRBN $T=850640 406680 0 0 $X=850640 $Y=406300
X1363 4855 718 4845 2 1 4871 QDFFRBN $T=851260 416760 1 0 $X=851260 $Y=411340
X1364 4870 4560 4768 2 1 4873 QDFFRBN $T=853740 487320 0 0 $X=853740 $Y=486940
X1365 4954 718 769 2 1 4908 QDFFRBN $T=872960 386520 0 180 $X=861180 $Y=381100
X1366 4912 718 4845 2 1 4939 QDFFRBN $T=861180 396600 0 0 $X=861180 $Y=396220
X1367 4913 696 4956 2 1 4949 QDFFRBN $T=861180 527640 1 0 $X=861180 $Y=522220
X1368 4960 4560 4935 2 1 4905 QDFFRBN $T=873580 467160 1 180 $X=861800 $Y=466780
X1369 4925 4560 4863 2 1 4948 QDFFRBN $T=863040 447000 1 0 $X=863040 $Y=441580
X1370 4927 4560 4935 2 1 4978 QDFFRBN $T=863040 487320 1 0 $X=863040 $Y=481900
X1371 4977 4560 4863 2 1 4929 QDFFRBN $T=875440 457080 1 180 $X=863660 $Y=456700
X1372 4931 4560 4956 2 1 4953 QDFFRBN $T=863660 507480 0 0 $X=863660 $Y=507100
X1373 4934 696 4956 2 1 780 QDFFRBN $T=863660 527640 0 0 $X=863660 $Y=527260
X1374 4924 4560 4768 2 1 4892 QDFFRBN $T=876060 497400 1 180 $X=864280 $Y=497020
X1375 4943 4560 4935 2 1 4952 QDFFRBN $T=865520 477240 1 0 $X=865520 $Y=471820
X1376 4973 718 4845 2 1 771 QDFFRBN $T=878540 416760 1 180 $X=866760 $Y=416380
X1377 5000 4560 4742 2 1 4950 QDFFRBN $T=883500 436920 1 180 $X=871720 $Y=436540
X1378 5022 4560 790 2 1 4976 QDFFRBN $T=884740 527640 0 180 $X=872960 $Y=522220
X1379 5036 718 769 2 1 4984 QDFFRBN $T=887220 386520 0 180 $X=875440 $Y=381100
X1380 4990 4560 5023 2 1 4993 QDFFRBN $T=876060 467160 0 0 $X=876060 $Y=466780
X1381 4991 4560 4935 2 1 5042 QDFFRBN $T=876060 487320 1 0 $X=876060 $Y=481900
X1382 807 696 796 2 1 782 QDFFRBN $T=887840 527640 1 180 $X=876060 $Y=527260
X1383 4997 4560 4863 2 1 4998 QDFFRBN $T=877300 457080 0 0 $X=877300 $Y=456700
X1384 5043 4560 4956 2 1 4995 QDFFRBN $T=889080 507480 1 180 $X=877300 $Y=507100
X1385 5026 4560 4742 2 1 4992 QDFFRBN $T=890940 436920 0 180 $X=879160 $Y=431500
X1386 5034 4560 4989 2 1 5003 QDFFRBN $T=890940 447000 0 180 $X=879160 $Y=441580
X1387 5011 718 769 2 1 802 QDFFRBN $T=879780 366360 0 0 $X=879780 $Y=365980
X1388 5047 718 4845 2 1 4987 QDFFRBN $T=892800 426840 0 180 $X=881020 $Y=421420
X1389 5076 4560 4956 2 1 5030 QDFFRBN $T=896520 507480 0 180 $X=884740 $Y=502060
X1390 5031 4560 4956 2 1 5085 QDFFRBN $T=884740 517560 0 0 $X=884740 $Y=517180
X1391 5075 718 769 2 1 793 QDFFRBN $T=897760 376440 1 180 $X=885980 $Y=376060
X1392 5028 718 4893 2 1 4999 QDFFRBN $T=898380 416760 0 180 $X=886600 $Y=411340
X1393 5055 4560 4989 2 1 5001 QDFFRBN $T=898380 436920 1 180 $X=886600 $Y=436540
X1394 5044 718 5081 2 1 5071 QDFFRBN $T=887220 406680 0 0 $X=887220 $Y=406300
X1395 5046 718 5081 2 1 5066 QDFFRBN $T=887840 396600 0 0 $X=887840 $Y=396220
X1396 5052 4560 4989 2 1 5102 QDFFRBN $T=889080 467160 1 0 $X=889080 $Y=461740
X1397 5056 4560 5023 2 1 5110 QDFFRBN $T=889700 467160 0 0 $X=889700 $Y=466780
X1398 5060 696 796 2 1 5097 QDFFRBN $T=890320 537720 1 0 $X=890320 $Y=532300
X1399 5061 4560 4989 2 1 814 QDFFRBN $T=890940 457080 0 0 $X=890940 $Y=456700
X1400 5062 696 790 2 1 5099 QDFFRBN $T=890940 527640 0 0 $X=890940 $Y=527260
X1401 5068 4560 4989 2 1 816 QDFFRBN $T=891560 447000 1 0 $X=891560 $Y=441580
X1402 5064 4560 4989 2 1 5123 QDFFRBN $T=891560 457080 1 0 $X=891560 $Y=451660
X1403 5065 4560 5098 2 1 795 QDFFRBN $T=891560 507480 0 0 $X=891560 $Y=507100
X1404 5059 718 809 2 1 4946 QDFFRBN $T=903960 376440 0 180 $X=892180 $Y=371020
X1405 5074 4560 4742 2 1 5087 QDFFRBN $T=892800 436920 1 0 $X=892800 $Y=431500
X1406 5079 718 4893 2 1 5113 QDFFRBN $T=894660 426840 1 0 $X=894660 $Y=421420
X1407 5129 820 5098 2 1 5078 QDFFRBN $T=907060 497400 0 180 $X=895280 $Y=491980
X1408 5156 820 5023 2 1 5080 QDFFRBN $T=907680 487320 0 180 $X=895900 $Y=481900
X1409 5094 718 809 2 1 5142 QDFFRBN $T=897140 366360 0 0 $X=897140 $Y=365980
X1410 5149 718 809 2 1 5093 QDFFRBN $T=908920 386520 0 180 $X=897140 $Y=381100
X1411 5106 4560 5158 2 1 5173 QDFFRBN $T=900860 436920 0 0 $X=900860 $Y=436540
X1412 5118 718 4893 2 1 812 QDFFRBN $T=913260 416760 0 180 $X=901480 $Y=411340
X1413 5124 820 5098 2 1 5141 QDFFRBN $T=903340 527640 1 0 $X=903340 $Y=522220
X1414 5183 718 5081 2 1 5112 QDFFRBN $T=916360 406680 0 180 $X=904580 $Y=401260
X1415 5131 820 5098 2 1 5190 QDFFRBN $T=904580 507480 1 0 $X=904580 $Y=502060
X1416 832 820 790 2 1 822 QDFFRBN $T=916360 537720 0 180 $X=904580 $Y=532300
X1417 5140 718 5158 2 1 5199 QDFFRBN $T=906440 406680 0 0 $X=906440 $Y=406300
X1418 5151 820 5098 2 1 5177 QDFFRBN $T=907060 497400 0 0 $X=907060 $Y=497020
X1419 5170 718 5081 2 1 5111 QDFFRBN $T=920080 386520 1 180 $X=908300 $Y=386140
X1420 5215 718 5081 2 1 826 QDFFRBN $T=920700 386520 0 180 $X=908920 $Y=381100
X1421 5159 718 5158 2 1 841 QDFFRBN $T=908920 426840 1 0 $X=908920 $Y=421420
X1422 5206 820 5023 2 1 5128 QDFFRBN $T=920700 467160 1 180 $X=908920 $Y=466780
X1423 5160 718 5158 2 1 5234 QDFFRBN $T=909540 436920 1 0 $X=909540 $Y=431500
X1424 5187 820 5023 2 1 5119 QDFFRBN $T=921320 487320 0 180 $X=909540 $Y=481900
X1425 5200 820 5184 2 1 5171 QDFFRBN $T=923180 457080 0 180 $X=911400 $Y=451660
X1426 5209 820 5158 2 1 5108 QDFFRBN $T=925040 447000 0 180 $X=913260 $Y=441580
X1427 5182 820 5098 2 1 5174 QDFFRBN $T=913880 517560 0 0 $X=913880 $Y=517180
X1428 5250 718 836 2 1 5198 QDFFRBN $T=929380 376440 1 180 $X=917600 $Y=376060
X1429 5216 820 5254 2 1 5139 QDFFRBN $T=920700 497400 0 0 $X=920700 $Y=497020
X1430 5217 820 849 2 1 5244 QDFFRBN $T=920700 527640 0 0 $X=920700 $Y=527260
X1431 5220 820 5184 2 1 858 QDFFRBN $T=921320 447000 0 0 $X=921320 $Y=446620
X1432 5268 718 5236 2 1 5211 QDFFRBN $T=933720 406680 0 180 $X=921940 $Y=401260
X1433 5228 820 5158 2 1 5260 QDFFRBN $T=921940 436920 0 0 $X=921940 $Y=436540
X1434 5223 820 5261 2 1 5267 QDFFRBN $T=921940 467160 1 0 $X=921940 $Y=461740
X1435 5218 846 5236 2 1 5230 QDFFRBN $T=922560 416760 0 0 $X=922560 $Y=416380
X1436 5208 820 5261 2 1 834 QDFFRBN $T=923180 477240 0 0 $X=923180 $Y=476860
X1437 5229 820 5254 2 1 5237 QDFFRBN $T=923180 487320 0 0 $X=923180 $Y=486940
X1438 847 718 859 2 1 854 QDFFRBN $T=925040 366360 0 0 $X=925040 $Y=365980
X1439 5294 846 836 2 1 5264 QDFFRBN $T=942400 376440 1 180 $X=930620 $Y=376060
X1440 5288 820 5266 2 1 853 QDFFRBN $T=944260 436920 0 180 $X=932480 $Y=431500
X1441 5276 846 5266 2 1 5311 QDFFRBN $T=933100 426840 1 0 $X=933100 $Y=421420
X1442 5317 820 5184 2 1 5274 QDFFRBN $T=944880 447000 1 180 $X=933100 $Y=446620
X1443 5325 820 5261 2 1 5280 QDFFRBN $T=946120 457080 1 180 $X=934340 $Y=456700
X1444 5319 846 5236 2 1 869 QDFFRBN $T=947360 406680 0 180 $X=935580 $Y=401260
X1445 5277 820 5261 2 1 856 QDFFRBN $T=947360 467160 0 180 $X=935580 $Y=461740
X1446 5287 820 5285 2 1 5296 QDFFRBN $T=935580 507480 0 0 $X=935580 $Y=507100
X1447 5293 820 5266 2 1 891 QDFFRBN $T=936820 436920 0 0 $X=936820 $Y=436540
X1448 5308 820 5254 2 1 5295 QDFFRBN $T=949220 487320 0 180 $X=937440 $Y=481900
X1449 5299 820 5254 2 1 5314 QDFFRBN $T=938060 477240 0 0 $X=938060 $Y=476860
X1450 5306 846 5236 2 1 878 QDFFRBN $T=952940 406680 1 180 $X=941160 $Y=406300
X1451 5330 846 883 2 1 5302 QDFFRBN $T=954180 376440 1 180 $X=942400 $Y=376060
X1452 5334 846 5364 2 1 5310 QDFFRBN $T=945500 416760 0 0 $X=945500 $Y=416380
X1453 5380 846 5328 2 1 5335 QDFFRBN $T=958520 416760 0 180 $X=946740 $Y=411340
X1454 5337 846 5364 2 1 898 QDFFRBN $T=946740 426840 1 0 $X=946740 $Y=421420
X1455 5336 820 5285 2 1 892 QDFFRBN $T=947360 507480 1 0 $X=947360 $Y=502060
X1456 5384 820 5285 2 1 5340 QDFFRBN $T=959140 517560 0 180 $X=947360 $Y=512140
X1457 5346 820 5285 2 1 5339 QDFFRBN $T=959140 527640 0 180 $X=947360 $Y=522220
X1458 5342 820 5376 2 1 5365 QDFFRBN $T=947980 467160 0 0 $X=947980 $Y=466780
X1459 5347 846 5379 2 1 901 QDFFRBN $T=948600 406680 1 0 $X=948600 $Y=401260
X1460 5373 820 5254 2 1 5343 QDFFRBN $T=961620 487320 0 180 $X=949840 $Y=481900
X1461 5355 820 918 2 1 887 QDFFRBN $T=950460 537720 1 0 $X=950460 $Y=532300
X1462 5386 820 5266 2 1 5361 QDFFRBN $T=964720 436920 1 180 $X=952940 $Y=436540
X1463 5414 846 5381 2 1 902 QDFFRBN $T=965960 376440 1 180 $X=954180 $Y=376060
X1464 5391 846 917 2 1 895 QDFFRBN $T=967200 376440 0 180 $X=955420 $Y=371020
X1465 5420 820 5348 2 1 5387 QDFFRBN $T=970300 447000 1 180 $X=958520 $Y=446620
X1466 5390 846 5364 2 1 5436 QDFFRBN $T=959140 416760 0 0 $X=959140 $Y=416380
X1467 5383 846 5379 2 1 5359 QDFFRBN $T=971540 386520 1 180 $X=959760 $Y=386140
X1468 5370 846 5266 2 1 910 QDFFRBN $T=972160 436920 0 180 $X=960380 $Y=431500
X1469 5426 820 5408 2 1 5395 QDFFRBN $T=972160 457080 1 180 $X=960380 $Y=456700
X1470 5417 820 5408 2 1 5389 QDFFRBN $T=972780 467160 1 180 $X=961000 $Y=466780
X1471 5400 820 5427 2 1 5374 QDFFRBN $T=961000 517560 1 0 $X=961000 $Y=512140
X1472 5398 820 918 2 1 872 QDFFRBN $T=972780 527640 0 180 $X=961000 $Y=522220
X1473 5394 846 5379 2 1 890 QDFFRBN $T=974020 396600 1 180 $X=962240 $Y=396220
X1474 5419 846 5379 2 1 886 QDFFRBN $T=974020 406680 0 180 $X=962240 $Y=401260
X1475 5411 846 5429 2 1 5448 QDFFRBN $T=963480 416760 1 0 $X=963480 $Y=411340
X1476 5428 820 5427 2 1 5392 QDFFRBN $T=975880 487320 0 180 $X=964100 $Y=481900
X1477 5409 820 5408 2 1 5377 QDFFRBN $T=975880 487320 1 180 $X=964100 $Y=486940
X1478 5397 820 5408 2 1 905 QDFFRBN $T=975880 497400 1 180 $X=964100 $Y=497020
X1479 5415 820 929 2 1 935 QDFFRBN $T=964720 537720 1 0 $X=964720 $Y=532300
X1480 5418 820 929 2 1 940 QDFFRBN $T=965340 517560 0 0 $X=965340 $Y=517180
X1481 5422 846 5381 2 1 938 QDFFRBN $T=965960 376440 0 0 $X=965960 $Y=376060
X1482 5423 820 5427 2 1 5441 QDFFRBN $T=965960 507480 1 0 $X=965960 $Y=502060
X1483 5432 846 5381 2 1 947 QDFFRBN $T=969060 386520 1 0 $X=969060 $Y=381100
X1484 5433 820 5456 2 1 5401 QDFFRBN $T=970300 447000 0 0 $X=970300 $Y=446620
X1485 950 846 926 2 1 903 QDFFRBN $T=982700 366360 1 180 $X=970920 $Y=365980
X1486 5476 846 5381 2 1 927 QDFFRBN $T=982700 376440 0 180 $X=970920 $Y=371020
X1487 5435 846 5328 2 1 5480 QDFFRBN $T=970920 406680 0 0 $X=970920 $Y=406300
X1488 5438 846 5429 2 1 5430 QDFFRBN $T=971540 426840 0 0 $X=971540 $Y=426460
X1489 5487 943 5376 2 1 5437 QDFFRBN $T=983320 477240 0 180 $X=971540 $Y=471820
X1490 5439 820 5456 2 1 945 QDFFRBN $T=974020 436920 0 0 $X=974020 $Y=436540
X1491 5458 943 5376 2 1 923 QDFFRBN $T=985800 467160 1 180 $X=974020 $Y=466780
X1492 5482 943 5427 2 1 5446 QDFFRBN $T=985800 517560 0 180 $X=974020 $Y=512140
X1493 5492 943 5456 2 1 5434 QDFFRBN $T=986420 457080 0 180 $X=974640 $Y=451660
X1494 5453 943 5427 2 1 5471 QDFFRBN $T=977120 497400 1 0 $X=977120 $Y=491980
X1495 941 943 929 2 1 967 QDFFRBN $T=977120 537720 1 0 $X=977120 $Y=532300
X1496 5469 943 5427 2 1 974 QDFFRBN $T=979600 477240 0 0 $X=979600 $Y=476860
X1497 5470 943 929 2 1 5532 QDFFRBN $T=979600 517560 0 0 $X=979600 $Y=517180
X1498 5473 943 929 2 1 977 QDFFRBN $T=980220 527640 1 0 $X=980220 $Y=522220
X1499 5485 820 5429 2 1 5525 QDFFRBN $T=983320 436920 1 0 $X=983320 $Y=431500
X1500 5505 846 926 2 1 5537 QDFFRBN $T=986420 366360 0 0 $X=986420 $Y=365980
X1501 5557 846 5328 2 1 5488 QDFFRBN $T=999440 416760 0 180 $X=987660 $Y=411340
X1502 5562 943 5456 2 1 5491 QDFFRBN $T=1000060 436920 1 180 $X=988280 $Y=436540
X1503 5513 943 5545 2 1 5524 QDFFRBN $T=988280 467160 0 0 $X=988280 $Y=466780
X1504 5572 943 5456 2 1 5523 QDFFRBN $T=1001920 457080 0 180 $X=990140 $Y=451660
X1505 5507 846 5547 2 1 5496 QDFFRBN $T=991380 386520 0 0 $X=991380 $Y=386140
X1506 5531 846 5547 2 1 972 QDFFRBN $T=1003160 396600 1 180 $X=991380 $Y=396220
X1507 5497 943 5456 2 1 5493 QDFFRBN $T=1003780 447000 1 180 $X=992000 $Y=446620
X1508 5536 943 5556 2 1 5528 QDFFRBN $T=992000 507480 1 0 $X=992000 $Y=502060
X1509 5539 943 5545 2 1 5551 QDFFRBN $T=992620 497400 1 0 $X=992620 $Y=491980
X1510 5542 846 5547 2 1 5553 QDFFRBN $T=993240 386520 1 0 $X=993240 $Y=381100
X1511 5544 943 5577 2 1 987 QDFFRBN $T=993240 517560 0 0 $X=993240 $Y=517180
X1512 5546 943 5556 2 1 5552 QDFFRBN $T=993860 517560 1 0 $X=993860 $Y=512140
X1513 5584 943 5556 2 1 5541 QDFFRBN $T=1006260 477240 1 180 $X=994480 $Y=476860
X1514 989 846 5547 2 1 1010 QDFFRBN $T=1000680 366360 0 0 $X=1000680 $Y=365980
X1515 5575 943 5628 2 1 5564 QDFFRBN $T=1000680 436920 0 0 $X=1000680 $Y=436540
X1516 1014 943 1000 2 1 988 QDFFRBN $T=1014940 537720 0 180 $X=1003160 $Y=532300
X1517 5635 846 5547 2 1 5606 QDFFRBN $T=1017420 386520 0 180 $X=1005640 $Y=381100
X1518 5598 943 5556 2 1 5663 QDFFRBN $T=1005640 497400 0 0 $X=1005640 $Y=497020
X1519 5620 943 5577 2 1 5609 QDFFRBN $T=1006880 517560 1 0 $X=1006880 $Y=512140
X1520 5629 846 5594 2 1 5587 QDFFRBN $T=1019280 396600 1 180 $X=1007500 $Y=396220
X1521 5665 943 5577 2 1 5624 QDFFRBN $T=1019280 527640 0 180 $X=1007500 $Y=522220
X1522 5619 943 5651 2 1 5610 QDFFRBN $T=1008120 467160 1 0 $X=1008120 $Y=461740
X1523 5622 943 5651 2 1 5602 QDFFRBN $T=1008120 467160 0 0 $X=1008120 $Y=466780
X1524 5654 846 5594 2 1 997 QDFFRBN $T=1020520 376440 0 180 $X=1008740 $Y=371020
X1525 5630 943 5651 2 1 1008 QDFFRBN $T=1008740 477240 1 0 $X=1008740 $Y=471820
X1526 5627 943 5348 2 1 5647 QDFFRBN $T=1009980 457080 1 0 $X=1009980 $Y=451660
X1527 5643 846 5628 2 1 5633 QDFFRBN $T=1023000 416760 0 180 $X=1011220 $Y=411340
X1528 5661 846 5628 2 1 5634 QDFFRBN $T=1023000 436920 0 180 $X=1011220 $Y=431500
X1529 5666 846 5628 2 1 5591 QDFFRBN $T=1023620 406680 0 180 $X=1011840 $Y=401260
X1530 5636 846 5628 2 1 5618 QDFFRBN $T=1023620 426840 0 180 $X=1011840 $Y=421420
X1531 5657 943 5651 2 1 5639 QDFFRBN $T=1024240 487320 0 180 $X=1012460 $Y=481900
X1532 5684 943 5577 2 1 1006 QDFFRBN $T=1024240 507480 0 180 $X=1012460 $Y=502060
X1533 1027 846 5547 2 1 1012 QDFFRBN $T=1026720 366360 1 180 $X=1014940 $Y=365980
X1534 5672 846 5628 2 1 5650 QDFFRBN $T=1026720 436920 1 180 $X=1014940 $Y=436540
X1535 5664 846 5594 2 1 5692 QDFFRBN $T=1016800 386520 0 0 $X=1016800 $Y=386140
X1536 1035 943 1000 2 1 1013 QDFFRBN $T=1028580 537720 0 180 $X=1016800 $Y=532300
X1537 5667 943 5690 2 1 1019 QDFFRBN $T=1018040 497400 0 0 $X=1018040 $Y=497020
X1538 5675 943 5690 2 1 5702 QDFFRBN $T=1020520 477240 0 0 $X=1020520 $Y=476860
X1539 5677 943 5651 2 1 5698 QDFFRBN $T=1021140 457080 0 0 $X=1021140 $Y=456700
X1540 5721 943 5674 2 1 5638 QDFFRBN $T=1032920 527640 0 180 $X=1021140 $Y=522220
X1541 5671 846 5713 2 1 5682 QDFFRBN $T=1021760 396600 0 0 $X=1021760 $Y=396220
X1542 5679 846 5713 2 1 5660 QDFFRBN $T=1022380 396600 1 0 $X=1022380 $Y=391180
X1543 5683 846 5723 2 1 5703 QDFFRBN $T=1023620 426840 1 0 $X=1023620 $Y=421420
X1544 5678 943 5651 2 1 5686 QDFFRBN $T=1023620 457080 1 0 $X=1023620 $Y=451660
X1545 5689 846 5727 2 1 1043 QDFFRBN $T=1024860 436920 1 0 $X=1024860 $Y=431500
X1546 5695 846 5723 2 1 5717 QDFFRBN $T=1025480 416760 0 0 $X=1025480 $Y=416380
X1547 5734 943 5690 2 1 5694 QDFFRBN $T=1038500 507480 0 180 $X=1026720 $Y=502060
X1548 5744 943 5674 2 1 5706 QDFFRBN $T=1041600 527640 1 180 $X=1029820 $Y=527260
X1549 5733 943 5690 2 1 5714 QDFFRBN $T=1044080 487320 0 180 $X=1032300 $Y=481900
X1550 5770 943 5690 2 1 1041 QDFFRBN $T=1044700 487320 1 180 $X=1032920 $Y=486940
X1551 5781 1039 5748 2 1 5735 QDFFRBN $T=1046560 467160 0 180 $X=1034780 $Y=461740
X1552 5763 943 5674 2 1 1034 QDFFRBN $T=1046560 517560 1 180 $X=1034780 $Y=517180
X1553 5779 1039 5713 2 1 5739 QDFFRBN $T=1047180 396600 1 180 $X=1035400 $Y=396220
X1554 5786 1039 5594 2 1 5719 QDFFRBN $T=1047800 386520 1 180 $X=1036020 $Y=386140
X1555 5743 943 5690 2 1 5791 QDFFRBN $T=1036020 477240 0 0 $X=1036020 $Y=476860
X1556 5783 1039 5748 2 1 5729 QDFFRBN $T=1048420 436920 1 180 $X=1036640 $Y=436540
X1557 5780 1039 5723 2 1 5740 QDFFRBN $T=1049040 416760 1 180 $X=1037260 $Y=416380
X1558 5750 1039 5723 2 1 5747 QDFFRBN $T=1037880 436920 1 0 $X=1037880 $Y=431500
X1559 5755 1039 5748 2 1 5772 QDFFRBN $T=1038500 457080 1 0 $X=1038500 $Y=451660
X1560 5758 1039 1056 2 1 5731 QDFFRBN $T=1052140 376440 0 180 $X=1040360 $Y=371020
X1561 5764 1039 5723 2 1 5828 QDFFRBN $T=1040360 416760 1 0 $X=1040360 $Y=411340
X1562 5766 943 5807 2 1 5736 QDFFRBN $T=1041600 507480 1 0 $X=1041600 $Y=502060
X1563 1068 1066 1057 2 1 1055 QDFFRBN $T=1054000 537720 0 180 $X=1042220 $Y=532300
X1564 5831 1066 5807 2 1 5793 QDFFRBN $T=1058340 507480 1 180 $X=1046560 $Y=507100
X1565 5817 1066 5788 2 1 5785 QDFFRBN $T=1058340 527640 0 180 $X=1046560 $Y=522220
X1566 5775 943 5807 2 1 5797 QDFFRBN $T=1047180 487320 0 0 $X=1047180 $Y=486940
X1567 5802 1039 5751 2 1 1078 QDFFRBN $T=1048420 376440 0 0 $X=1048420 $Y=376060
X1568 5803 1039 5751 2 1 5850 QDFFRBN $T=1048420 386520 1 0 $X=1048420 $Y=381100
X1569 5808 1039 5751 2 1 5841 QDFFRBN $T=1049660 386520 0 0 $X=1049660 $Y=386140
X1570 5809 1039 5834 2 1 5801 QDFFRBN $T=1049660 396600 0 0 $X=1049660 $Y=396220
X1571 5812 1039 5727 2 1 5844 QDFFRBN $T=1050900 436920 0 0 $X=1050900 $Y=436540
X1572 5814 1039 5727 2 1 5826 QDFFRBN $T=1052140 436920 1 0 $X=1052140 $Y=431500
X1573 5866 1039 5834 2 1 5818 QDFFRBN $T=1064540 416760 1 180 $X=1052760 $Y=416380
X1574 5815 1039 5845 2 1 1060 QDFFRBN $T=1052760 457080 1 0 $X=1052760 $Y=451660
X1575 5821 1066 5845 2 1 5752 QDFFRBN $T=1052760 487320 1 0 $X=1052760 $Y=481900
X1576 5825 1066 5845 2 1 5813 QDFFRBN $T=1053380 477240 0 0 $X=1053380 $Y=476860
X1577 5876 1066 5845 2 1 1071 QDFFRBN $T=1067020 467160 0 180 $X=1055240 $Y=461740
X1578 5872 1039 5848 2 1 5835 QDFFRBN $T=1067640 447000 0 180 $X=1055860 $Y=441580
X1579 5863 1066 5807 2 1 5833 QDFFRBN $T=1067640 497400 1 180 $X=1055860 $Y=497020
X1580 5840 1066 5788 2 1 5820 QDFFRBN $T=1057100 517560 1 0 $X=1057100 $Y=512140
X1581 5908 1039 5834 2 1 5860 QDFFRBN $T=1073220 396600 1 180 $X=1061440 $Y=396220
X1582 5861 1066 5848 2 1 1074 QDFFRBN $T=1073220 457080 1 180 $X=1061440 $Y=456700
X1583 5851 1066 5807 2 1 5868 QDFFRBN $T=1061440 487320 0 0 $X=1061440 $Y=486940
X1584 5865 1066 5788 2 1 5885 QDFFRBN $T=1062680 527640 0 0 $X=1062680 $Y=527260
X1585 5922 1039 1056 2 1 5869 QDFFRBN $T=1076320 376440 0 180 $X=1064540 $Y=371020
X1586 5926 1039 5834 2 1 5874 QDFFRBN $T=1076940 416760 1 180 $X=1065160 $Y=416380
X1587 5887 1066 5845 2 1 5928 QDFFRBN $T=1067020 467160 1 0 $X=1067020 $Y=461740
X1588 5932 1039 5848 2 1 5890 QDFFRBN $T=1079420 436920 0 180 $X=1067640 $Y=431500
X1589 5930 1039 5848 2 1 5899 QDFFRBN $T=1080660 447000 0 180 $X=1068880 $Y=441580
X1590 5903 1066 5807 2 1 5917 QDFFRBN $T=1070120 497400 0 0 $X=1070120 $Y=497020
X1591 5939 1066 5788 2 1 5909 QDFFRBN $T=1083140 517560 1 180 $X=1071360 $Y=517180
X1592 5912 1039 5950 2 1 5889 QDFFRBN $T=1073220 426840 1 0 $X=1073220 $Y=421420
X1593 5915 1066 5951 2 1 5958 QDFFRBN $T=1073220 487320 1 0 $X=1073220 $Y=481900
X1594 5919 1039 5957 2 1 5941 QDFFRBN $T=1074460 386520 1 0 $X=1074460 $Y=381100
X1595 5949 1039 5913 2 1 5920 QDFFRBN $T=1086240 396600 1 180 $X=1074460 $Y=396220
X1596 5927 1039 5951 2 1 5937 QDFFRBN $T=1075080 457080 0 0 $X=1075080 $Y=456700
X1597 5921 1066 1100 2 1 5901 QDFFRBN $T=1075080 517560 1 0 $X=1075080 $Y=512140
X1598 5934 1066 5788 2 1 5960 QDFFRBN $T=1076320 527640 0 0 $X=1076320 $Y=527260
X1599 5936 1066 5951 2 1 5956 QDFFRBN $T=1076940 477240 0 0 $X=1076940 $Y=476860
X1600 5938 1039 5950 2 1 5968 QDFFRBN $T=1077560 436920 0 0 $X=1077560 $Y=436540
X1601 5947 1066 1100 2 1 6009 QDFFRBN $T=1080660 507480 1 0 $X=1080660 $Y=502060
X1602 6007 1039 5957 2 1 1094 QDFFRBN $T=1094300 366360 1 180 $X=1082520 $Y=365980
X1603 5965 1039 5957 2 1 1108 QDFFRBN $T=1083760 376440 1 0 $X=1083760 $Y=371020
X1604 5980 1066 5951 2 1 6021 QDFFRBN $T=1086860 487320 1 0 $X=1086860 $Y=481900
X1605 5977 1039 5990 2 1 5955 QDFFRBN $T=1087480 426840 1 0 $X=1087480 $Y=421420
X1606 5985 1039 6011 2 1 1110 QDFFRBN $T=1088100 457080 0 0 $X=1088100 $Y=456700
X1607 6037 1039 5913 2 1 5986 QDFFRBN $T=1100500 386520 1 180 $X=1088720 $Y=386140
X1608 5987 1066 5951 2 1 6018 QDFFRBN $T=1088720 487320 0 0 $X=1088720 $Y=486940
X1609 6032 1039 5990 2 1 5992 QDFFRBN $T=1101740 436920 0 180 $X=1089960 $Y=431500
X1610 6029 1039 6011 2 1 5972 QDFFRBN $T=1102360 447000 0 180 $X=1090580 $Y=441580
X1611 5998 1066 1114 2 1 5979 QDFFRBN $T=1091820 517560 1 0 $X=1091820 $Y=512140
X1612 6026 1039 5913 2 1 5995 QDFFRBN $T=1105460 396600 1 180 $X=1093680 $Y=396220
X1613 6057 1039 6011 2 1 6012 QDFFRBN $T=1105460 457080 0 180 $X=1093680 $Y=451660
X1614 6014 1066 1114 2 1 6016 QDFFRBN $T=1094300 507480 0 0 $X=1094300 $Y=507100
X1615 6047 1039 6033 2 1 5991 QDFFRBN $T=1106700 416760 0 180 $X=1094920 $Y=411340
X1616 6023 1039 5957 2 1 6059 QDFFRBN $T=1095540 376440 0 0 $X=1095540 $Y=376060
X1617 6051 1039 6011 2 1 6020 QDFFRBN $T=1107320 467160 0 180 $X=1095540 $Y=461740
X1618 6017 1066 1114 2 1 6041 QDFFRBN $T=1096780 527640 1 0 $X=1096780 $Y=522220
X1619 6071 1039 5950 2 1 6038 QDFFRBN $T=1111040 436920 1 180 $X=1099260 $Y=436540
X1620 6061 1066 5951 2 1 6030 QDFFRBN $T=1112280 487320 0 180 $X=1100500 $Y=481900
X1621 6094 1039 5913 2 1 6046 QDFFRBN $T=1112900 396600 0 180 $X=1101120 $Y=391180
X1622 6044 1039 6033 2 1 6008 QDFFRBN $T=1112900 426840 0 180 $X=1101120 $Y=421420
X1623 6103 1039 5913 2 1 6054 QDFFRBN $T=1114760 386520 1 180 $X=1102980 $Y=386140
X1624 6091 1039 6011 2 1 6045 QDFFRBN $T=1114760 457080 1 180 $X=1102980 $Y=456700
X1625 6062 1066 1114 2 1 6084 QDFFRBN $T=1104840 517560 1 0 $X=1104840 $Y=512140
X1626 6119 1066 1121 2 1 6056 QDFFRBN $T=1116620 537720 0 180 $X=1104840 $Y=532300
X1627 6081 1039 6033 2 1 6108 QDFFRBN $T=1108560 416760 1 0 $X=1108560 $Y=411340
X1628 6124 1039 5990 2 1 6105 QDFFRBN $T=1126540 436920 1 180 $X=1114760 $Y=436540
X1629 6136 1039 1126 2 1 6069 QDFFRBN $T=1127780 396600 0 180 $X=1116000 $Y=391180
X1630 6134 1039 6033 2 1 6095 QDFFRBN $T=1127780 426840 0 180 $X=1116000 $Y=421420
X1631 6089 1039 1126 2 1 1120 QDFFRBN $T=1128400 376440 0 180 $X=1116620 $Y=371020
X1632 6118 1039 1126 2 1 6036 QDFFRBN $T=1128400 376440 1 180 $X=1116620 $Y=376060
X1633 6123 1039 1126 2 1 6013 QDFFRBN $T=1128400 386520 1 180 $X=1116620 $Y=386140
X1634 6131 1039 1126 2 1 1119 QDFFRBN $T=1128400 406680 1 180 $X=1116620 $Y=406300
X1635 6140 1039 6033 2 1 6078 QDFFRBN $T=1128400 426840 1 180 $X=1116620 $Y=426460
X1636 6130 1066 6125 2 1 6088 QDFFRBN $T=1128400 457080 1 180 $X=1116620 $Y=456700
X1637 6129 1066 6125 2 1 6087 QDFFRBN $T=1128400 467160 0 180 $X=1116620 $Y=461740
X1638 6112 1066 6125 2 1 1117 QDFFRBN $T=1128400 467160 1 180 $X=1116620 $Y=466780
X1639 6116 1066 6125 2 1 6079 QDFFRBN $T=1128400 477240 1 180 $X=1116620 $Y=476860
X1640 6114 1066 6125 2 1 6082 QDFFRBN $T=1128400 487320 0 180 $X=1116620 $Y=481900
X1641 6117 1066 6138 2 1 6085 QDFFRBN $T=1116620 487320 0 0 $X=1116620 $Y=486940
X1642 6115 1066 6138 2 1 6076 QDFFRBN $T=1116620 497400 0 0 $X=1116620 $Y=497020
X1643 6127 1066 6138 2 1 6064 QDFFRBN $T=1116620 507480 1 0 $X=1116620 $Y=502060
X1644 6139 1039 6125 2 1 6102 QDFFRBN $T=1129020 447000 0 180 $X=1117240 $Y=441580
X1645 6126 1066 6138 2 1 6063 QDFFRBN $T=1117240 517560 1 0 $X=1117240 $Y=512140
X1646 6098 1066 1121 2 1 5774 QDFFRBN $T=1117240 517560 0 0 $X=1117240 $Y=517180
X1647 6128 1066 1121 2 1 6109 QDFFRBN $T=1117240 527640 0 0 $X=1117240 $Y=527260
X1648 2835 1 2 2831 2806 2774 1202 ICV_4 $T=500340 477240 0 0 $X=500340 $Y=476860
X1649 3551 1 2 3584 3587 3621 1202 ICV_4 $T=598300 527640 1 0 $X=598300 $Y=522220
X1650 3695 1 2 3735 3739 3758 1202 ICV_4 $T=620000 497400 0 0 $X=620000 $Y=497020
X1651 3784 1 2 3809 3811 3838 1202 ICV_4 $T=633640 497400 0 0 $X=633640 $Y=497020
X1652 3801 1 2 3820 3825 3851 1202 ICV_4 $T=636120 467160 1 0 $X=636120 $Y=461740
X1653 491 1 2 3842 3844 3872 1202 ICV_4 $T=639220 527640 1 0 $X=639220 $Y=522220
X1654 3857 1 2 3907 507 516 1202 ICV_4 $T=649760 457080 0 0 $X=649760 $Y=456700
X1655 3954 1 2 3973 3980 3992 1202 ICV_4 $T=661540 457080 1 0 $X=661540 $Y=451660
X1656 3956 1 2 3974 3983 3982 1202 ICV_4 $T=661540 517560 0 0 $X=661540 $Y=517180
X1657 3970 1 2 3987 3988 4003 1202 ICV_4 $T=663400 467160 0 0 $X=663400 $Y=466780
X1658 4012 1 2 4041 4046 4058 1202 ICV_4 $T=674560 537720 1 0 $X=674560 $Y=532300
X1659 3993 1 2 4027 4015 4045 1202 ICV_4 $T=677660 477240 1 0 $X=677660 $Y=471820
X1660 4052 1 2 4068 4072 4090 1202 ICV_4 $T=680140 426840 0 0 $X=680140 $Y=426460
X1661 4113 1 2 4132 4143 4163 1202 ICV_4 $T=692540 366360 0 0 $X=692540 $Y=365980
X1662 4144 1 2 4166 4137 4181 1202 ICV_4 $T=701220 477240 0 0 $X=701220 $Y=476860
X1663 4176 1 2 4168 4133 4153 1202 ICV_4 $T=705560 416760 1 0 $X=705560 $Y=411340
X1664 4098 1 2 4127 4209 4178 1202 ICV_4 $T=707420 507480 0 0 $X=707420 $Y=507100
X1665 4177 1 2 4225 4227 4248 1202 ICV_4 $T=716100 416760 1 0 $X=716100 $Y=411340
X1666 4224 1 2 4238 4221 4256 1202 ICV_4 $T=717960 376440 0 0 $X=717960 $Y=376060
X1667 4270 1 2 4304 4309 4332 1202 ICV_4 $T=727260 487320 1 0 $X=727260 $Y=481900
X1668 4280 1 2 4307 4312 4319 1202 ICV_4 $T=727880 457080 0 0 $X=727880 $Y=456700
X1669 4300 1 2 4297 4296 4292 1202 ICV_4 $T=734080 507480 1 0 $X=734080 $Y=502060
X1670 4447 1 2 4470 4473 4482 1202 ICV_4 $T=762600 487320 1 0 $X=762600 $Y=481900
X1671 4548 1 2 4564 4567 4575 1202 ICV_4 $T=783060 517560 0 0 $X=783060 $Y=517180
X1672 4556 1 2 4566 4571 4572 1202 ICV_4 $T=784300 457080 1 0 $X=784300 $Y=451660
X1673 4601 1 2 4604 4476 4544 1202 ICV_4 $T=796080 386520 1 0 $X=796080 $Y=381100
X1674 4569 1 2 4623 4602 4668 1202 ICV_4 $T=798560 376440 1 0 $X=798560 $Y=371020
X1675 4643 1 2 4630 4698 4701 1202 ICV_4 $T=811580 507480 0 0 $X=811580 $Y=507100
X1676 4645 1 2 4634 4673 4664 1202 ICV_4 $T=812200 487320 1 0 $X=812200 $Y=481900
X1677 4691 1 2 4708 690 4721 1202 ICV_4 $T=812820 376440 0 0 $X=812820 $Y=376060
X1678 4663 1 2 4678 4640 4639 1202 ICV_4 $T=812820 457080 0 0 $X=812820 $Y=456700
X1679 4744 1 2 4761 4738 4759 1202 ICV_4 $T=828320 517560 1 0 $X=828320 $Y=512140
X1680 4816 1 2 4811 4835 4829 1202 ICV_4 $T=842580 416760 0 0 $X=842580 $Y=416380
X1681 4769 1 2 4777 743 4879 1202 ICV_4 $T=846300 537720 1 0 $X=846300 $Y=532300
X1682 4871 1 2 4885 4900 4919 1202 ICV_4 $T=854360 416760 0 0 $X=854360 $Y=416380
X1683 4873 1 2 4896 4892 4897 1202 ICV_4 $T=854360 497400 1 0 $X=854360 $Y=491980
X1684 4949 1 2 4972 4978 4965 1202 ICV_4 $T=871720 497400 1 0 $X=871720 $Y=491980
X1685 4976 1 2 4996 4681 4589 1202 ICV_4 $T=879780 537720 1 0 $X=879780 $Y=532300
X1686 5003 1 2 5017 4993 5020 1202 ICV_4 $T=881020 457080 1 0 $X=881020 $Y=451660
X1687 4992 1 2 5013 4999 5004 1202 ICV_4 $T=884120 416760 0 0 $X=884120 $Y=416380
X1688 5030 1 2 5049 5035 5058 1202 ICV_4 $T=884740 497400 0 0 $X=884740 $Y=497020
X1689 4939 1 2 4967 5066 5067 1202 ICV_4 $T=887220 386520 1 0 $X=887220 $Y=381100
X1690 5001 1 2 5039 4948 4975 1202 ICV_4 $T=890940 447000 0 0 $X=890940 $Y=446620
X1691 5087 1 2 5095 5113 5114 1202 ICV_4 $T=897140 416760 0 0 $X=897140 $Y=416380
X1692 5099 1 2 5103 5097 5086 1202 ICV_4 $T=902720 527640 0 0 $X=902720 $Y=527260
X1693 4995 1 2 5024 5296 5329 1202 ICV_4 $T=962240 497400 1 0 $X=962240 $Y=491980
X1694 5190 1 2 5176 5257 5197 1202 ICV_4 $T=962240 527640 0 0 $X=962240 $Y=527260
X1695 5395 1 2 5431 5434 5445 1202 ICV_4 $T=964720 467160 1 0 $X=964720 $Y=461740
X1696 5387 1 2 5407 5401 5425 1202 ICV_4 $T=970300 447000 1 0 $X=970300 $Y=441580
X1697 5491 1 2 5514 5493 5526 1202 ICV_4 $T=984560 447000 1 0 $X=984560 $Y=441580
X1698 5537 1 2 5540 5553 5559 1202 ICV_4 $T=992620 376440 0 0 $X=992620 $Y=376060
X1699 5609 1 2 5632 5638 5653 1202 ICV_4 $T=1005640 517560 0 0 $X=1005640 $Y=517180
X1700 5610 1 2 5608 5647 5637 1202 ICV_4 $T=1008740 457080 0 0 $X=1008740 $Y=456700
X1701 5591 1 2 5646 5634 5649 1202 ICV_4 $T=1013700 416760 0 0 $X=1013700 $Y=416380
X1702 1022 1 2 1031 5698 5697 1202 ICV_4 $T=1021140 487320 0 0 $X=1021140 $Y=486940
X1703 5650 1 2 5659 5714 5711 1202 ICV_4 $T=1024860 467160 1 0 $X=1024860 $Y=461740
X1704 5717 1 2 5722 5740 5759 1202 ICV_4 $T=1030440 416760 1 0 $X=1030440 $Y=411340
X1705 5729 1 2 5745 5735 5769 1202 ICV_4 $T=1032920 457080 0 0 $X=1032920 $Y=456700
X1706 5901 1 2 5914 5917 5916 1202 ICV_4 $T=1068880 507480 1 0 $X=1068880 $Y=502060
X1707 5899 1 2 5910 5972 5993 1202 ICV_4 $T=1080660 447000 1 0 $X=1080660 $Y=441580
X1708 5968 1 2 5978 5992 6001 1202 ICV_4 $T=1086240 426840 0 0 $X=1086240 $Y=426460
X1709 1106 1 2 1112 1113 1116 1202 ICV_4 $T=1092440 537720 1 0 $X=1092440 $Y=532300
X1710 5991 1 2 6031 5995 6010 1202 ICV_4 $T=1097400 406680 1 0 $X=1097400 $Y=401260
X1711 6036 1 2 6055 6059 6060 1202 ICV_4 $T=1099260 376440 1 0 $X=1099260 $Y=371020
X1712 5833 1 2 5882 6012 6083 1202 ICV_4 $T=1101740 436920 1 0 $X=1101740 $Y=431500
X1713 6082 1 2 6092 6079 6096 1202 ICV_4 $T=1115380 477240 1 0 $X=1115380 $Y=471820
X1714 6102 1 2 6132 6087 6100 1202 ICV_4 $T=1119720 457080 1 0 $X=1119720 $Y=451660
X1715 6063 1 2 6107 6084 6110 1202 ICV_4 $T=1119720 507480 0 0 $X=1119720 $Y=507100
X1716 1321 1243 2 1 44 1331 MUX2 $T=243040 527640 1 0 $X=243040 $Y=522220
X1717 1777 1758 2 1 1735 1766 MUX2 $T=320540 467160 1 180 $X=316200 $Y=466780
X1718 1773 1758 2 1 1809 1790 MUX2 $T=318060 416760 1 0 $X=318060 $Y=411340
X1719 1753 1758 2 1 1762 1799 MUX2 $T=318060 436920 0 0 $X=318060 $Y=436540
X1720 1763 1758 2 1 1782 1776 MUX2 $T=318060 457080 1 0 $X=318060 $Y=451660
X1721 1676 112 2 1 1779 1806 MUX2 $T=318680 376440 1 0 $X=318680 $Y=371020
X1722 1771 1785 2 1 1792 1812 MUX2 $T=320540 386520 0 0 $X=320540 $Y=386140
X1723 1772 1785 2 1 1813 1807 MUX2 $T=320540 406680 1 0 $X=320540 $Y=401260
X1724 1760 1785 2 1 1827 1816 MUX2 $T=321780 406680 0 0 $X=321780 $Y=406300
X1725 1786 1795 2 1 1754 1820 MUX2 $T=321780 477240 0 0 $X=321780 $Y=476860
X1726 1742 1785 2 1 1810 1764 MUX2 $T=323020 376440 0 0 $X=323020 $Y=376060
X1727 1804 1758 2 1 1793 1836 MUX2 $T=325500 426840 1 0 $X=325500 $Y=421420
X1728 1811 1785 2 1 1859 1822 MUX2 $T=327360 396600 1 0 $X=327360 $Y=391180
X1729 1843 1795 2 1 1842 1869 MUX2 $T=332940 487320 0 0 $X=332940 $Y=486940
X1730 1890 1795 2 1 1846 1866 MUX2 $T=341620 487320 1 180 $X=337280 $Y=486940
X1731 2239 2408 2 1 2394 2390 MUX2 $T=426560 467160 1 180 $X=422220 $Y=466780
X1732 2290 2408 2 1 2439 2422 MUX2 $T=424700 467160 1 0 $X=424700 $Y=461740
X1733 2073 2408 2 1 2441 2442 MUX2 $T=426560 467160 0 0 $X=426560 $Y=466780
X1734 2461 1795 2 1 2436 2410 MUX2 $T=434620 487320 0 180 $X=430280 $Y=481900
X1735 2472 2408 2 1 2494 2489 MUX2 $T=435860 467160 0 0 $X=435860 $Y=466780
X1736 2491 2457 2 1 2483 2484 MUX2 $T=442060 487320 1 180 $X=437720 $Y=486940
X1737 2527 2457 2 1 2506 2462 MUX2 $T=445160 497400 1 180 $X=440820 $Y=497020
X1738 252 249 2 1 2508 2507 MUX2 $T=445160 517560 0 180 $X=440820 $Y=512140
X1739 2543 249 2 1 2553 2564 MUX2 $T=446400 517560 0 0 $X=446400 $Y=517180
X1740 2634 2631 2 1 2538 2549 MUX2 $T=463140 507480 0 180 $X=458800 $Y=502060
X1741 269 2631 2 1 2654 2629 MUX2 $T=461900 507480 0 0 $X=461900 $Y=507100
X1742 2623 2631 2 1 2663 2682 MUX2 $T=463760 507480 1 0 $X=463760 $Y=502060
X1743 2741 2748 2 1 2728 2774 MUX2 $T=481120 477240 0 0 $X=481120 $Y=476860
X1744 299 295 2 1 2768 2790 MUX2 $T=483600 507480 0 0 $X=483600 $Y=507100
X1745 2781 2811 2 1 2740 2782 MUX2 $T=491660 457080 0 180 $X=487320 $Y=451660
X1746 2804 2748 2 1 2767 2831 MUX2 $T=490420 477240 0 0 $X=490420 $Y=476860
X1747 2785 2811 2 1 2766 2754 MUX2 $T=492280 457080 1 0 $X=492280 $Y=451660
X1748 2818 2811 2 1 2765 2845 MUX2 $T=492900 447000 0 0 $X=492900 $Y=446620
X1749 2850 2811 2 1 2873 2872 MUX2 $T=497240 467160 1 0 $X=497240 $Y=461740
X1750 2848 295 2 1 2868 326 MUX2 $T=504060 527640 1 180 $X=499720 $Y=527260
X1751 2917 295 2 1 2807 2886 MUX2 $T=507780 517560 0 180 $X=503440 $Y=512140
X1752 355 2948 2 1 3082 3033 MUX2 $T=522040 396600 0 0 $X=522040 $Y=396220
X1753 3176 3117 2 1 3076 346 MUX2 $T=534440 517560 0 180 $X=530100 $Y=512140
X1754 3148 3117 2 1 3166 374 MUX2 $T=533200 507480 0 0 $X=533200 $Y=507100
X1755 3126 3191 2 1 3148 3054 MUX2 $T=540640 507480 0 180 $X=536300 $Y=502060
X1756 3095 3191 2 1 3176 372 MUX2 $T=541880 507480 1 180 $X=537540 $Y=507100
X1757 3268 3117 2 1 3219 391 MUX2 $T=551180 507480 1 180 $X=546840 $Y=507100
X1758 3222 2948 2 1 3124 3243 MUX2 $T=553040 406680 1 180 $X=548700 $Y=406300
X1759 3271 3117 2 1 3214 401 MUX2 $T=551180 507480 0 0 $X=551180 $Y=507100
X1760 3303 3296 2 1 2978 397 MUX2 $T=556760 376440 1 180 $X=552420 $Y=376060
X1761 3284 399 2 1 3252 3313 MUX2 $T=553660 386520 0 0 $X=553660 $Y=386140
X1762 3108 3296 2 1 3225 3334 MUX2 $T=554280 376440 1 0 $X=554280 $Y=371020
X1763 3284 3180 2 1 3158 3318 MUX2 $T=554280 406680 1 0 $X=554280 $Y=401260
X1764 3292 3191 2 1 3270 3322 MUX2 $T=555520 426840 1 0 $X=555520 $Y=421420
X1765 405 3191 2 1 3268 3095 MUX2 $T=559860 507480 1 180 $X=555520 $Y=507100
X1766 3326 3296 2 1 3186 3303 MUX2 $T=561100 376440 1 180 $X=556760 $Y=376060
X1767 3340 3296 2 1 392 404 MUX2 $T=562960 366360 1 180 $X=558620 $Y=365980
X1768 3326 399 2 1 2997 3304 MUX2 $T=562960 396600 0 180 $X=558620 $Y=391180
X1769 3318 3296 2 1 3237 3272 MUX2 $T=562960 406680 0 180 $X=558620 $Y=401260
X1770 3025 3191 2 1 3224 2982 MUX2 $T=564200 497400 0 180 $X=559860 $Y=491980
X1771 407 3191 2 1 3271 405 MUX2 $T=564200 507480 0 180 $X=559860 $Y=502060
X1772 3966 3967 2 1 3918 517 MUX2 $T=663400 497400 1 180 $X=659060 $Y=497020
X1773 3982 523 2 1 3935 3963 MUX2 $T=667120 517560 0 180 $X=662780 $Y=512140
X1774 3991 3967 2 1 3945 520 MUX2 $T=668980 527640 1 180 $X=664640 $Y=527260
X1775 3974 3967 2 1 3936 3963 MUX2 $T=671460 517560 0 180 $X=667120 $Y=512140
X1776 3996 523 2 1 3989 517 MUX2 $T=672700 487320 1 180 $X=668360 $Y=486940
X1777 4027 4022 2 1 3944 520 MUX2 $T=676420 467160 0 180 $X=672080 $Y=461740
X1778 4003 4036 2 1 3957 520 MUX2 $T=677660 467160 1 180 $X=673320 $Y=466780
X1779 4045 4036 2 1 3943 517 MUX2 $T=680140 457080 1 180 $X=675800 $Y=456700
X1780 4058 4053 2 1 3998 3963 MUX2 $T=680140 517560 0 180 $X=675800 $Y=512140
X1781 3973 4022 2 1 4030 4070 MUX2 $T=680760 457080 1 0 $X=680760 $Y=451660
X1782 4091 4036 2 1 4065 4070 MUX2 $T=689440 457080 1 180 $X=685100 $Y=456700
X1783 4114 4105 2 1 4040 4070 MUX2 $T=693780 436920 0 180 $X=689440 $Y=431500
X1784 4128 4119 2 1 4042 548 MUX2 $T=695640 467160 1 180 $X=691300 $Y=466780
X1785 4171 4120 2 1 4110 548 MUX2 $T=699360 517560 1 180 $X=695020 $Y=517180
X1786 4187 4089 2 1 4147 4070 MUX2 $T=706800 436920 0 180 $X=702460 $Y=431500
X1787 4166 4099 2 1 4189 548 MUX2 $T=702460 477240 1 0 $X=702460 $Y=471820
X1788 4132 4172 2 1 4169 4070 MUX2 $T=708040 376440 1 180 $X=703700 $Y=376060
X1789 4090 4105 2 1 4232 4240 MUX2 $T=714240 447000 1 0 $X=714240 $Y=441580
X1790 579 4215 2 1 583 4070 MUX2 $T=714860 376440 1 0 $X=714860 $Y=371020
X1791 4218 4197 2 1 4236 4228 MUX2 $T=714860 497400 1 0 $X=714860 $Y=491980
X1792 4225 4089 2 1 4241 4245 MUX2 $T=716720 426840 1 0 $X=716720 $Y=421420
X1793 585 4173 2 1 4190 4228 MUX2 $T=722300 527640 1 180 $X=717960 $Y=527260
X1794 4230 4231 2 1 4257 4245 MUX2 $T=719200 416760 0 0 $X=719200 $Y=416380
X1795 4238 4215 2 1 4266 4245 MUX2 $T=719820 376440 1 0 $X=719820 $Y=371020
X1796 4269 4220 2 1 4246 4240 MUX2 $T=725400 447000 1 180 $X=721060 $Y=446620
X1797 4248 4239 2 1 4273 4245 MUX2 $T=721680 396600 0 0 $X=721680 $Y=396220
X1798 4249 564 2 1 4275 4228 MUX2 $T=721680 507480 1 0 $X=721680 $Y=502060
X1799 4256 4172 2 1 4278 4245 MUX2 $T=722920 386520 0 0 $X=722920 $Y=386140
X1800 4274 4188 2 1 4261 4255 MUX2 $T=730360 477240 0 180 $X=726020 $Y=471820
X1801 4297 4276 2 1 4244 4228 MUX2 $T=730980 517560 1 180 $X=726640 $Y=517180
X1802 4319 4324 2 1 4279 4245 MUX2 $T=734080 447000 0 180 $X=729740 $Y=441580
X1803 4308 4205 2 1 4318 4315 MUX2 $T=732220 467160 0 0 $X=732220 $Y=466780
X1804 592 582 2 1 4234 599 MUX2 $T=732220 537720 1 0 $X=732220 $Y=532300
X1805 4321 4173 2 1 4334 599 MUX2 $T=734080 527640 1 0 $X=734080 $Y=522220
X1806 4331 4205 2 1 4345 4255 MUX2 $T=736560 467160 0 0 $X=736560 $Y=466780
X1807 3759 4276 2 1 4311 4351 MUX2 $T=737800 517560 1 0 $X=737800 $Y=512140
X1808 4358 4210 2 1 4337 4339 MUX2 $T=743380 436920 0 180 $X=739040 $Y=431500
X1809 4341 4215 2 1 4350 4359 MUX2 $T=739660 376440 0 0 $X=739660 $Y=376060
X1810 4357 4268 2 1 4342 4339 MUX2 $T=744000 426840 0 180 $X=739660 $Y=421420
X1811 4343 3995 2 1 4366 4351 MUX2 $T=740280 497400 0 0 $X=740280 $Y=497020
X1812 4307 4348 2 1 4361 4315 MUX2 $T=740900 467160 0 0 $X=740900 $Y=466780
X1813 608 4322 2 1 4277 4359 MUX2 $T=741520 386520 1 0 $X=741520 $Y=381100
X1814 4370 4324 2 1 4340 4339 MUX2 $T=747100 447000 0 180 $X=742760 $Y=441580
X1815 617 4231 2 1 4333 4339 MUX2 $T=748340 426840 0 180 $X=744000 $Y=421420
X1816 4381 4382 2 1 4362 4351 MUX2 $T=748960 487320 1 180 $X=744620 $Y=486940
X1817 620 564 2 1 611 613 MUX2 $T=748960 537720 0 180 $X=744620 $Y=532300
X1818 4393 4220 2 1 4413 4339 MUX2 $T=751440 457080 1 0 $X=751440 $Y=451660
X1819 4304 4400 2 1 4355 613 MUX2 $T=755780 517560 1 180 $X=751440 $Y=517180
X1820 4396 4356 2 1 4346 4414 MUX2 $T=752060 386520 0 0 $X=752060 $Y=386140
X1821 3899 4400 2 1 4397 4399 MUX2 $T=756400 487320 1 180 $X=752060 $Y=486940
X1822 4405 4401 2 1 4421 4407 MUX2 $T=753300 406680 0 0 $X=753300 $Y=406300
X1823 633 4239 2 1 4378 4407 MUX2 $T=758260 416760 1 180 $X=753920 $Y=416380
X1824 4411 4356 2 1 4417 4429 MUX2 $T=755160 376440 0 0 $X=755160 $Y=376060
X1825 3668 4382 2 1 4432 634 MUX2 $T=755780 527640 1 0 $X=755780 $Y=522220
X1826 3693 4400 2 1 4435 4436 MUX2 $T=757020 487320 0 0 $X=757020 $Y=486940
X1827 3924 4400 2 1 4375 4423 MUX2 $T=761360 517560 1 180 $X=757020 $Y=517180
X1828 3987 4416 2 1 4445 4399 MUX2 $T=759500 467160 0 0 $X=759500 $Y=466780
X1829 4001 4385 2 1 4454 4407 MUX2 $T=760120 447000 1 0 $X=760120 $Y=441580
X1830 636 4400 2 1 4469 634 MUX2 $T=760120 527640 1 0 $X=760120 $Y=522220
X1831 3758 4400 2 1 4386 4464 MUX2 $T=761360 507480 1 0 $X=761360 $Y=502060
X1832 4452 4401 2 1 4451 4414 MUX2 $T=763840 386520 0 0 $X=763840 $Y=386140
X1833 4478 4444 2 1 4428 4407 MUX2 $T=768180 426840 1 180 $X=763840 $Y=426460
X1834 4470 4426 2 1 4455 4399 MUX2 $T=768180 467160 1 180 $X=763840 $Y=466780
X1835 4482 4382 2 1 4458 4464 MUX2 $T=770040 497400 1 180 $X=765700 $Y=497020
X1836 4491 4401 2 1 4427 4429 MUX2 $T=770660 376440 1 180 $X=766320 $Y=376060
X1837 4487 4382 2 1 4442 4423 MUX2 $T=770660 517560 0 180 $X=766320 $Y=512140
X1838 4474 4382 2 1 4493 4436 MUX2 $T=767560 487320 0 0 $X=767560 $Y=486940
X1839 3584 629 2 1 4495 4496 MUX2 $T=775620 527640 1 180 $X=771280 $Y=527260
X1840 3951 4416 2 1 4522 4459 MUX2 $T=772520 467160 0 0 $X=772520 $Y=466780
X1841 4335 4444 2 1 4488 4507 MUX2 $T=777480 426840 0 180 $X=773140 $Y=421420
X1842 4510 4239 2 1 4468 649 MUX2 $T=773760 406680 0 0 $X=773760 $Y=406300
X1843 4463 4415 2 1 4500 649 MUX2 $T=781200 447000 0 180 $X=776860 $Y=441580
X1844 3809 4513 2 1 4526 4399 MUX2 $T=781200 497400 0 180 $X=776860 $Y=491980
X1845 4437 4524 2 1 4552 4459 MUX2 $T=776860 497400 0 0 $X=776860 $Y=497020
X1846 4529 4430 2 1 4545 4507 MUX2 $T=778100 416760 0 0 $X=778100 $Y=416380
X1847 4534 4401 2 1 4547 649 MUX2 $T=778720 406680 0 0 $X=778720 $Y=406300
X1848 4538 4356 2 1 4561 656 MUX2 $T=779960 396600 0 0 $X=779960 $Y=396220
X1849 4540 4385 2 1 4549 4507 MUX2 $T=780580 436920 0 0 $X=780580 $Y=436540
X1850 4544 4401 2 1 4532 656 MUX2 $T=781820 386520 0 0 $X=781820 $Y=386140
X1851 4554 4401 2 1 4576 4550 MUX2 $T=784300 376440 0 0 $X=784300 $Y=376060
X1852 4551 4415 2 1 4559 4518 MUX2 $T=789260 436920 0 180 $X=784920 $Y=431500
X1853 4574 4444 2 1 4543 4518 MUX2 $T=789880 406680 1 180 $X=785540 $Y=406300
X1854 4572 4416 2 1 4536 4464 MUX2 $T=789880 467160 1 180 $X=785540 $Y=466780
X1855 4566 4385 2 1 4558 4518 MUX2 $T=791740 436920 1 180 $X=787400 $Y=436540
X1856 4588 4426 2 1 4553 4464 MUX2 $T=794840 467160 1 180 $X=790500 $Y=466780
X1857 4564 629 2 1 4615 662 MUX2 $T=791120 527640 1 0 $X=791120 $Y=522220
X1858 4604 627 2 1 4565 4550 MUX2 $T=796700 376440 1 180 $X=792360 $Y=376060
X1859 4589 654 2 1 4613 4423 MUX2 $T=794220 527640 0 0 $X=794220 $Y=527260
X1860 664 4444 2 1 4619 4610 MUX2 $T=795460 416760 0 0 $X=795460 $Y=416380
X1861 666 4444 2 1 4629 4597 MUX2 $T=796700 406680 0 0 $X=796700 $Y=406300
X1862 4605 4415 2 1 4609 4610 MUX2 $T=801660 436920 1 180 $X=797320 $Y=436540
X1863 4625 4426 2 1 4595 4611 MUX2 $T=801660 477240 0 180 $X=797320 $Y=471820
X1864 4630 4513 2 1 4600 662 MUX2 $T=802280 507480 1 180 $X=797940 $Y=507100
X1865 4634 4513 2 1 4585 4436 MUX2 $T=802900 487320 1 180 $X=798560 $Y=486940
X1866 4638 4415 2 1 4608 656 MUX2 $T=804140 447000 1 180 $X=799800 $Y=446620
X1867 4639 4416 2 1 4594 4617 MUX2 $T=804140 467160 1 180 $X=799800 $Y=466780
X1868 4623 627 2 1 4618 4429 MUX2 $T=801040 366360 0 0 $X=801040 $Y=365980
X1869 671 654 2 1 4647 680 MUX2 $T=801040 527640 0 0 $X=801040 $Y=527260
X1870 678 615 2 1 4627 4550 MUX2 $T=806620 376440 1 180 $X=802280 $Y=376060
X1871 674 4513 2 1 4665 4666 MUX2 $T=804140 487320 0 0 $X=804140 $Y=486940
X1872 4658 4415 2 1 4677 4682 MUX2 $T=806620 436920 0 0 $X=806620 $Y=436540
X1873 3872 4513 2 1 4689 4423 MUX2 $T=807240 507480 0 0 $X=807240 $Y=507100
X1874 4664 4416 2 1 4684 4610 MUX2 $T=807860 477240 0 0 $X=807860 $Y=476860
X1875 4668 615 2 1 4686 4429 MUX2 $T=808480 376440 1 0 $X=808480 $Y=371020
X1876 682 4426 2 1 4687 4610 MUX2 $T=808480 457080 0 0 $X=808480 $Y=456700
X1877 4671 4426 2 1 4688 4682 MUX2 $T=808480 467160 1 0 $X=808480 $Y=461740
X1878 683 4385 2 1 4692 656 MUX2 $T=809100 447000 0 0 $X=809100 $Y=446620
X1879 4662 4444 2 1 4696 4682 MUX2 $T=809720 406680 0 0 $X=809720 $Y=406300
X1880 4676 4385 2 1 4699 4682 MUX2 $T=810340 436920 1 0 $X=810340 $Y=431500
X1881 4678 4416 2 1 4706 4682 MUX2 $T=810340 467160 0 0 $X=810340 $Y=466780
X1882 4693 4524 2 1 4715 688 MUX2 $T=812820 507480 1 0 $X=812820 $Y=502060
X1883 687 4430 2 1 4711 4631 MUX2 $T=814680 406680 1 0 $X=814680 $Y=401260
X1884 4041 629 2 1 4720 680 MUX2 $T=815300 527640 1 0 $X=815300 $Y=522220
X1885 4708 4728 2 1 4680 4550 MUX2 $T=823360 386520 1 180 $X=819020 $Y=386140
X1886 693 4430 2 1 4716 4695 MUX2 $T=819020 406680 1 0 $X=819020 $Y=401260
X1887 4721 4725 2 1 695 4429 MUX2 $T=823980 366360 1 180 $X=819640 $Y=365980
X1888 4736 4728 2 1 4703 4429 MUX2 $T=827080 376440 1 180 $X=822740 $Y=376060
X1889 699 4728 2 1 697 637 MUX2 $T=828320 366360 1 180 $X=823980 $Y=365980
X1890 4749 4728 2 1 4723 4597 MUX2 $T=830180 406680 0 180 $X=825840 $Y=401260
X1891 4753 4739 2 1 4700 4737 MUX2 $T=830800 477240 0 180 $X=826460 $Y=471820
X1892 4741 4728 2 1 4747 684 MUX2 $T=827080 376440 0 0 $X=827080 $Y=376060
X1893 700 4725 2 1 712 637 MUX2 $T=828320 366360 0 0 $X=828320 $Y=365980
X1894 4764 4725 2 1 4718 4597 MUX2 $T=834520 406680 0 180 $X=830180 $Y=401260
X1895 4775 4725 2 1 4727 684 MUX2 $T=835760 386520 0 180 $X=831420 $Y=381100
X1896 4782 4781 2 1 4760 705 MUX2 $T=836380 507480 0 180 $X=832040 $Y=502060
X1897 4759 4739 2 1 4792 705 MUX2 $T=833280 497400 0 0 $X=833280 $Y=497020
X1898 4771 4725 2 1 4788 4737 MUX2 $T=834520 406680 1 0 $X=834520 $Y=401260
X1899 4777 711 2 1 4802 721 MUX2 $T=835140 537720 1 0 $X=835140 $Y=532300
X1900 730 732 2 1 723 722 MUX2 $T=843820 537720 0 180 $X=839480 $Y=532300
X1901 724 4725 2 1 4731 4631 MUX2 $T=840100 386520 0 0 $X=840100 $Y=386140
X1902 734 4822 2 1 4745 4812 MUX2 $T=846300 517560 0 180 $X=841960 $Y=512140
X1903 4829 4820 2 1 4798 4812 MUX2 $T=846920 497400 1 180 $X=842580 $Y=497020
X1904 4831 4828 2 1 728 729 MUX2 $T=847540 366360 1 180 $X=843200 $Y=365980
X1905 4821 4820 2 1 4840 4255 MUX2 $T=843820 467160 1 0 $X=843820 $Y=461740
X1906 4838 4828 2 1 4824 4631 MUX2 $T=849400 386520 1 180 $X=845060 $Y=386140
X1907 4761 4820 2 1 4807 731 MUX2 $T=850020 487320 1 180 $X=845680 $Y=486940
X1908 4832 4830 2 1 4850 4737 MUX2 $T=846920 406680 1 0 $X=846920 $Y=401260
X1909 742 4849 2 1 738 729 MUX2 $T=851880 366360 1 180 $X=847540 $Y=365980
X1910 4856 4822 2 1 4826 4255 MUX2 $T=851880 467160 1 180 $X=847540 $Y=466780
X1911 4878 4876 2 1 4837 4812 MUX2 $T=855600 507480 1 180 $X=851260 $Y=507100
X1912 753 4849 2 1 4813 745 MUX2 $T=856220 366360 1 180 $X=851880 $Y=365980
X1913 4885 4883 2 1 4855 745 MUX2 $T=858080 406680 0 180 $X=853740 $Y=401260
X1914 762 4898 2 1 4810 4812 MUX2 $T=859320 517560 1 180 $X=854980 $Y=517180
X1915 754 4828 2 1 764 745 MUX2 $T=856220 366360 0 0 $X=856220 $Y=365980
X1916 4896 4876 2 1 4870 756 MUX2 $T=860560 487320 0 180 $X=856220 $Y=481900
X1917 4884 4886 2 1 4904 4732 MUX2 $T=856840 426840 0 0 $X=856840 $Y=426460
X1918 758 759 2 1 4890 722 MUX2 $T=856840 527640 0 0 $X=856840 $Y=527260
X1919 4906 4886 2 1 4842 4631 MUX2 $T=861800 396600 0 180 $X=857460 $Y=391180
X1920 4919 4922 2 1 4851 745 MUX2 $T=862420 406680 0 180 $X=858080 $Y=401260
X1921 4920 4923 2 1 4888 4732 MUX2 $T=863040 436920 0 180 $X=858700 $Y=431500
X1922 4938 4883 2 1 4954 729 MUX2 $T=865520 386520 0 0 $X=865520 $Y=386140
X1923 4961 4964 2 1 4931 4812 MUX2 $T=870480 507480 0 180 $X=866140 $Y=502060
X1924 4944 4926 2 1 4960 4917 MUX2 $T=866760 467160 1 0 $X=866760 $Y=461740
X1925 4967 4922 2 1 4912 729 MUX2 $T=871720 396600 0 180 $X=867380 $Y=391180
X1926 4963 4958 2 1 4945 4631 MUX2 $T=871720 406680 1 180 $X=867380 $Y=406300
X1927 4969 4971 2 1 4943 756 MUX2 $T=871720 477240 1 180 $X=867380 $Y=476860
X1928 4965 4964 2 1 4927 756 MUX2 $T=871720 497400 0 180 $X=867380 $Y=491980
X1929 4972 4971 2 1 4913 4812 MUX2 $T=871720 517560 1 180 $X=867380 $Y=517180
X1930 781 4951 2 1 787 784 MUX2 $T=871100 376440 1 0 $X=871100 $Y=371020
X1931 788 783 2 1 5011 797 MUX2 $T=876060 376440 1 0 $X=876060 $Y=371020
X1932 4996 4971 2 1 5022 806 MUX2 $T=877920 517560 0 0 $X=877920 $Y=517180
X1933 5020 4964 2 1 4990 4917 MUX2 $T=883500 467160 0 180 $X=879160 $Y=461740
X1934 5004 4883 2 1 5028 5038 MUX2 $T=879780 406680 0 0 $X=879780 $Y=406300
X1935 5013 5014 2 1 5026 4732 MUX2 $T=880400 426840 0 0 $X=880400 $Y=426460
X1936 5017 4971 2 1 5034 4732 MUX2 $T=881640 447000 0 0 $X=881640 $Y=446620
X1937 5018 800 2 1 5036 5038 MUX2 $T=882880 386520 0 0 $X=882880 $Y=386140
X1938 5041 4971 2 1 4997 4917 MUX2 $T=887840 467160 0 180 $X=883500 $Y=461740
X1939 5024 5027 2 1 5043 5038 MUX2 $T=883500 497400 1 0 $X=883500 $Y=491980
X1940 5006 5033 2 1 5047 4732 MUX2 $T=884740 426840 0 0 $X=884740 $Y=426460
X1941 5039 4964 2 1 5055 4732 MUX2 $T=886600 447000 0 0 $X=886600 $Y=446620
X1942 5063 4739 2 1 4991 5037 MUX2 $T=892180 487320 0 180 $X=887840 $Y=481900
X1943 5067 4922 2 1 5046 797 MUX2 $T=892800 396600 0 180 $X=888460 $Y=391180
X1944 5049 4781 2 1 5076 5038 MUX2 $T=888460 497400 1 0 $X=888460 $Y=491980
X1945 5053 808 2 1 5075 5038 MUX2 $T=889700 386520 0 0 $X=889700 $Y=386140
X1946 5077 5083 2 1 5031 5037 MUX2 $T=894660 517560 0 180 $X=890320 $Y=512140
X1947 5086 5083 2 1 5060 806 MUX2 $T=896520 527640 0 180 $X=892180 $Y=522220
X1948 5103 4841 2 1 5062 806 MUX2 $T=900860 527640 0 180 $X=896520 $Y=522220
X1949 815 4964 2 1 5065 5038 MUX2 $T=902100 497400 1 180 $X=897760 $Y=497020
X1950 811 4922 2 1 5118 4695 MUX2 $T=899000 406680 1 0 $X=899000 $Y=401260
X1951 5120 5027 2 1 5056 5096 MUX2 $T=903340 477240 1 180 $X=899000 $Y=476860
X1952 5105 5082 2 1 5129 821 MUX2 $T=900860 487320 0 0 $X=900860 $Y=486940
X1953 5117 5122 2 1 5149 784 MUX2 $T=902720 386520 0 0 $X=902720 $Y=386140
X1954 5134 5027 2 1 5156 821 MUX2 $T=905200 487320 0 0 $X=905200 $Y=486940
X1955 5148 4922 2 1 5170 784 MUX2 $T=907680 396600 1 0 $X=907680 $Y=391180
X1956 5175 4841 2 1 5124 5045 MUX2 $T=912640 517560 1 180 $X=908300 $Y=517180
X1957 5176 5126 2 1 5131 821 MUX2 $T=913260 517560 0 180 $X=908920 $Y=512140
X1958 5178 5126 2 1 5151 5096 MUX2 $T=913880 497400 0 180 $X=909540 $Y=491980
X1959 5180 4951 2 1 5094 827 MUX2 $T=914500 376440 0 180 $X=910160 $Y=371020
X1960 5166 5122 2 1 5183 827 MUX2 $T=910780 396600 0 0 $X=910780 $Y=396220
X1961 835 5192 2 1 5208 5207 MUX2 $T=915740 477240 1 0 $X=915740 $Y=471820
X1962 5197 4915 2 1 5224 5179 MUX2 $T=918840 527640 1 0 $X=918840 $Y=522220
X1963 5205 5122 2 1 5140 833 MUX2 $T=919460 406680 0 0 $X=919460 $Y=406300
X1964 848 4876 2 1 5225 5207 MUX2 $T=926900 477240 0 180 $X=922560 $Y=471820
X1965 5255 5259 2 1 5217 5179 MUX2 $T=928140 527640 0 180 $X=923800 $Y=522220
X1966 5243 5212 2 1 5268 5240 MUX2 $T=926900 406680 0 0 $X=926900 $Y=406300
X1967 5248 5104 2 1 5252 5249 MUX2 $T=933720 507480 1 180 $X=929380 $Y=507100
X1968 5315 4915 2 1 5282 5045 MUX2 $T=939300 527640 0 180 $X=934960 $Y=522220
X1969 5318 5104 2 1 5299 5207 MUX2 $T=942400 477240 0 180 $X=938060 $Y=471820
X1970 5324 5321 2 1 5308 5207 MUX2 $T=944260 487320 1 180 $X=939920 $Y=486940
X1971 5329 5048 2 1 5287 5249 MUX2 $T=946120 507480 0 180 $X=941780 $Y=502060
X1972 5360 5104 2 1 5346 5045 MUX2 $T=952940 517560 1 180 $X=948600 $Y=517180
X1973 900 5338 2 1 5370 904 MUX2 $T=951080 436920 1 0 $X=951080 $Y=431500
X1974 911 5048 2 1 5355 5045 MUX2 $T=957280 517560 1 180 $X=952940 $Y=517180
X1975 5371 5332 2 1 5386 904 MUX2 $T=954800 447000 1 0 $X=954800 $Y=441580
X1976 913 5259 2 1 5398 5410 MUX2 $T=957280 517560 0 0 $X=957280 $Y=517180
X1977 5404 5321 2 1 5384 5249 MUX2 $T=962240 507480 1 180 $X=957900 $Y=507100
X1978 920 912 2 1 5414 904 MUX2 $T=961620 366360 0 0 $X=961620 $Y=365980
X1979 5424 5259 2 1 5400 5249 MUX2 $T=967200 507480 1 180 $X=962860 $Y=507100
X1980 5445 5466 2 1 5492 956 MUX2 $T=979600 457080 0 0 $X=979600 $Y=456700
X1981 5502 5442 2 1 5435 5240 MUX2 $T=985180 416760 0 180 $X=980840 $Y=411340
X1982 5526 5457 2 1 5497 956 MUX2 $T=990140 447000 1 180 $X=985800 $Y=446620
X1983 5540 942 2 1 5505 904 MUX2 $T=993860 376440 0 180 $X=989520 $Y=371020
X1984 5530 5444 2 1 5557 5240 MUX2 $T=991380 416760 0 0 $X=991380 $Y=416380
X1985 5646 5571 2 1 5666 5554 MUX2 $T=1013700 406680 0 0 $X=1013700 $Y=406300
X1986 5656 5640 2 1 5679 5668 MUX2 $T=1016180 396600 1 0 $X=1016180 $Y=391180
X1987 5685 5596 2 1 5671 5668 MUX2 $T=1024860 406680 1 180 $X=1020520 $Y=406300
X1988 5691 5596 2 1 5664 5554 MUX2 $T=1026100 376440 1 180 $X=1021760 $Y=376060
X1989 5701 5527 2 1 5675 1023 MUX2 $T=1026100 477240 0 180 $X=1021760 $Y=471820
X1990 5705 5615 2 1 5683 1023 MUX2 $T=1029200 426840 1 180 $X=1024860 $Y=426460
X1991 5711 5699 2 1 5733 1023 MUX2 $T=1030440 477240 1 0 $X=1030440 $Y=471820
X1992 5741 980 2 1 5758 5554 MUX2 $T=1036020 376440 0 0 $X=1036020 $Y=376060
X1993 5759 5603 2 1 5780 5668 MUX2 $T=1039740 406680 0 0 $X=1039740 $Y=406300
X1994 5777 5771 2 1 5743 5765 MUX2 $T=1045320 477240 0 180 $X=1040980 $Y=471820
X1995 5756 5762 2 1 5766 5765 MUX2 $T=1045320 507480 1 180 $X=1040980 $Y=507100
X1996 5738 1042 2 1 5786 5668 MUX2 $T=1042840 386520 1 0 $X=1042840 $Y=381100
X1997 5795 5642 2 1 5775 5765 MUX2 $T=1047800 497400 0 180 $X=1043460 $Y=491980
X1998 5794 5789 2 1 5809 1063 MUX2 $T=1047180 406680 1 0 $X=1047180 $Y=401260
X1999 5799 5644 2 1 5817 1067 MUX2 $T=1048420 517560 0 0 $X=1048420 $Y=517180
X2000 5822 1061 2 1 1062 1063 MUX2 $T=1054000 366360 1 180 $X=1049660 $Y=365980
X2001 5811 5687 2 1 5831 1067 MUX2 $T=1050280 517560 1 0 $X=1050280 $Y=512140
X2002 5839 5790 2 1 5764 1065 MUX2 $T=1056480 406680 1 180 $X=1052140 $Y=406300
X2003 5849 5699 2 1 5825 5765 MUX2 $T=1059580 477240 0 180 $X=1055240 $Y=471820
X2004 5867 5842 2 1 5851 5847 MUX2 $T=1063920 497400 0 180 $X=1059580 $Y=491980
X2005 5855 5854 2 1 5866 1065 MUX2 $T=1060820 426840 1 0 $X=1060820 $Y=421420
X2006 5879 5790 2 1 5837 5859 MUX2 $T=1066400 406680 1 180 $X=1062060 $Y=406300
X2007 5882 5858 2 1 5863 5859 MUX2 $T=1067020 507480 1 180 $X=1062680 $Y=507100
X2008 5883 5852 2 1 5865 5859 MUX2 $T=1067020 527640 0 180 $X=1062680 $Y=522220
X2009 5806 5810 2 1 5894 5895 MUX2 $T=1064540 426840 0 0 $X=1064540 $Y=426460
X2010 5888 5789 2 1 5908 5895 MUX2 $T=1067640 406680 0 0 $X=1067640 $Y=406300
X2011 5902 1083 2 1 5922 5856 MUX2 $T=1069500 376440 0 0 $X=1069500 $Y=376060
X2012 1089 5881 2 1 5876 5847 MUX2 $T=1069500 477240 1 0 $X=1069500 $Y=471820
X2013 1090 1061 2 1 1092 5856 MUX2 $T=1070120 366360 0 0 $X=1070120 $Y=365980
X2014 5773 5900 2 1 5821 5847 MUX2 $T=1070120 477240 0 0 $X=1070120 $Y=476860
X2015 5906 5790 2 1 5919 5918 MUX2 $T=1070740 396600 1 0 $X=1070740 $Y=391180
X2016 5904 5905 2 1 5932 5847 MUX2 $T=1070740 436920 0 0 $X=1070740 $Y=436540
X2017 5864 5852 2 1 5878 5907 MUX2 $T=1075080 527640 0 180 $X=1070740 $Y=522220
X2018 5910 5880 2 1 5930 5847 MUX2 $T=1071980 457080 1 0 $X=1071980 $Y=451660
X2019 5931 5900 2 1 5887 5911 MUX2 $T=1076320 467160 1 180 $X=1071980 $Y=466780
X2020 5914 5858 2 1 5921 5410 MUX2 $T=1078800 507480 1 180 $X=1074460 $Y=507100
X2021 5952 1042 2 1 5923 5918 MUX2 $T=1079420 366360 1 180 $X=1075080 $Y=365980
X2022 5924 5836 2 1 5939 5907 MUX2 $T=1075080 527640 1 0 $X=1075080 $Y=522220
X2023 5929 5789 2 1 5926 5859 MUX2 $T=1076320 406680 0 0 $X=1076320 $Y=406300
X2024 5935 5789 2 1 5949 5918 MUX2 $T=1076940 406680 1 0 $X=1076940 $Y=401260
X2025 5945 5880 2 1 5927 5895 MUX2 $T=1081280 457080 0 180 $X=1076940 $Y=451660
X2026 5946 5842 2 1 5915 5911 MUX2 $T=1081280 487320 1 180 $X=1076940 $Y=486940
X2027 5959 5881 2 1 5936 5911 MUX2 $T=1083140 467160 1 180 $X=1078800 $Y=466780
X2028 5974 5836 2 1 5934 1093 MUX2 $T=1083760 527640 0 180 $X=1079420 $Y=522220
X2029 5978 5905 2 1 5938 5895 MUX2 $T=1086860 447000 1 180 $X=1082520 $Y=446620
X2030 6002 5789 2 1 5953 5969 MUX2 $T=1089960 406680 1 180 $X=1085620 $Y=406300
X2031 1107 5900 2 1 5985 5907 MUX2 $T=1093680 477240 0 180 $X=1089340 $Y=471820
X2032 6004 5852 2 1 5998 5999 MUX2 $T=1094920 517560 1 180 $X=1090580 $Y=517180
X2033 6001 5905 2 1 6032 5969 MUX2 $T=1091200 436920 0 0 $X=1091200 $Y=436540
X2034 6015 5881 2 1 5980 1103 MUX2 $T=1095540 477240 1 180 $X=1091200 $Y=476860
X2035 6022 5842 2 1 5987 6003 MUX2 $T=1096160 497400 1 180 $X=1091820 $Y=497020
X2036 6006 5790 2 1 6037 6027 MUX2 $T=1092440 396600 1 0 $X=1092440 $Y=391180
X2037 6024 5852 2 1 5996 1093 MUX2 $T=1096780 527640 0 180 $X=1092440 $Y=522220
X2038 6010 5789 2 1 6026 6027 MUX2 $T=1093060 406680 0 0 $X=1093060 $Y=406300
X2039 5993 5880 2 1 6029 5969 MUX2 $T=1093060 447000 0 0 $X=1093060 $Y=446620
X2040 6040 5858 2 1 6014 6003 MUX2 $T=1100500 497400 1 180 $X=1096160 $Y=497020
X2041 1109 1061 2 1 6007 6043 MUX2 $T=1096780 366360 0 0 $X=1096780 $Y=365980
X2042 6028 5810 2 1 6044 1115 MUX2 $T=1096780 416760 0 0 $X=1096780 $Y=416380
X2043 6031 5790 2 1 6047 1115 MUX2 $T=1097400 406680 0 0 $X=1097400 $Y=406300
X2044 6060 1084 2 1 6023 1115 MUX2 $T=1105460 366360 1 180 $X=1101120 $Y=365980
X2045 6048 5900 2 1 6061 1103 MUX2 $T=1101120 477240 0 0 $X=1101120 $Y=476860
X2046 6083 5880 2 1 6057 5918 MUX2 $T=1109180 447000 1 180 $X=1104840 $Y=446620
X2047 6101 5905 2 1 6071 5918 MUX2 $T=1111040 447000 0 180 $X=1106700 $Y=441580
X2048 6110 5858 2 1 6062 6074 MUX2 $T=1111660 507480 1 180 $X=1107320 $Y=507100
X2049 6055 1084 2 1 6118 6043 MUX2 $T=1109180 376440 1 0 $X=1109180 $Y=371020
X2050 6111 5854 2 1 6081 6043 MUX2 $T=1113520 406680 1 180 $X=1109180 $Y=406300
X2051 1122 5900 2 1 6112 1123 MUX2 $T=1109180 467160 1 0 $X=1109180 $Y=461740
X2052 6113 1083 2 1 6089 1115 MUX2 $T=1114760 366360 1 180 $X=1110420 $Y=365980
X2053 6092 5881 2 1 6114 6074 MUX2 $T=1110420 477240 0 0 $X=1110420 $Y=476860
X2054 6086 5858 2 1 6127 6099 MUX2 $T=1110420 507480 1 0 $X=1110420 $Y=502060
X2055 6090 5810 2 1 6094 6043 MUX2 $T=1115380 396600 1 180 $X=1111040 $Y=396220
X2056 6096 5900 2 1 6116 6074 MUX2 $T=1111040 477240 1 0 $X=1111040 $Y=471820
X2057 6097 5842 2 1 6117 6074 MUX2 $T=1111040 487320 0 0 $X=1111040 $Y=486940
X2058 6104 1083 2 1 6123 6027 MUX2 $T=1112280 386520 1 0 $X=1112280 $Y=381100
X2059 6106 5905 2 1 6124 1123 MUX2 $T=1112280 447000 1 0 $X=1112280 $Y=441580
X2060 6107 5852 2 1 6126 6099 MUX2 $T=1112280 517560 0 0 $X=1112280 $Y=517180
X2061 6120 5905 2 1 6130 6074 MUX2 $T=1115380 447000 0 0 $X=1115380 $Y=446620
X2062 6121 5836 2 1 6119 6080 MUX2 $T=1115380 527640 1 0 $X=1115380 $Y=522220
X2063 1125 5854 2 1 6131 6027 MUX2 $T=1116000 396600 0 0 $X=1116000 $Y=396220
X2064 6122 5854 2 1 6134 1095 MUX2 $T=1116000 416760 0 0 $X=1116000 $Y=416380
X2065 6132 5880 2 1 6139 1123 MUX2 $T=1119720 447000 0 0 $X=1119720 $Y=446620
X2066 6137 5852 2 1 6128 6080 MUX2 $T=1124060 527640 0 180 $X=1119720 $Y=522220
X2067 6133 5810 2 1 6136 6027 MUX2 $T=1120340 396600 0 0 $X=1120340 $Y=396220
X2068 6135 5810 2 1 6140 1095 MUX2 $T=1121580 416760 0 0 $X=1121580 $Y=416380
X2069 139 1922 1941 1942 1 145 2 AOI22S $T=350920 376440 0 0 $X=350920 $Y=376060
X2070 1840 139 1952 143 1 1960 2 AOI22S $T=355260 386520 0 180 $X=351540 $Y=381100
X2071 2855 2834 2793 2827 1 2788 2 AOI22S $T=497860 426840 0 180 $X=494140 $Y=421420
X2072 2952 343 2959 344 1 2984 2 AOI22S $T=512120 376440 1 0 $X=512120 $Y=371020
X2073 2894 350 3012 3015 1 2984 2 AOI22S $T=517080 386520 1 0 $X=517080 $Y=381100
X2074 3014 350 3013 3026 1 354 2 AOI22S $T=517700 376440 0 0 $X=517700 $Y=376060
X2075 2953 354 3022 3015 1 2984 2 AOI22S $T=518320 386520 0 0 $X=518320 $Y=386140
X2076 3076 2771 3096 2584 1 3048 2 AOI22S $T=525760 487320 1 180 $X=522040 $Y=486940
X2077 3102 370 3097 3015 1 2984 2 AOI22S $T=528860 386520 1 180 $X=525140 $Y=386140
X2078 3014 366 3071 3026 1 371 2 AOI22S $T=525140 396600 1 0 $X=525140 $Y=391180
X2079 3056 367 3079 2993 1 3045 2 AOI22S $T=525140 416760 0 0 $X=525140 $Y=416380
X2080 3014 369 3059 3026 1 373 2 AOI22S $T=525760 376440 0 0 $X=525760 $Y=376060
X2081 3114 366 3109 3015 1 2984 2 AOI22S $T=530100 386520 0 180 $X=526380 $Y=381100
X2082 3014 359 3036 3026 1 352 2 AOI22S $T=526380 396600 0 0 $X=526380 $Y=396220
X2083 3100 369 379 344 1 360 2 AOI22S $T=533200 366360 1 180 $X=529480 $Y=365980
X2084 3111 352 3121 2993 1 3045 2 AOI22S $T=529480 416760 0 0 $X=529480 $Y=416380
X2085 2843 376 3144 3015 1 3045 2 AOI22S $T=532580 386520 1 0 $X=532580 $Y=381100
X2086 3025 3150 3127 3148 1 3107 2 AOI22S $T=532580 507480 1 0 $X=532580 $Y=502060
X2087 3153 371 3170 3015 1 3045 2 AOI22S $T=536920 386520 1 180 $X=533200 $Y=386140
X2088 3174 359 3169 2993 1 3045 2 AOI22S $T=537540 416760 1 180 $X=533820 $Y=416380
X2089 3166 3150 3184 3025 1 3205 2 AOI22S $T=538160 497400 0 0 $X=538160 $Y=497020
X2090 3198 355 3206 383 1 3033 2 AOI22S $T=540640 396600 1 0 $X=540640 $Y=391180
X2091 3223 3161 3217 3204 1 3134 2 AOI22S $T=544360 487320 0 180 $X=540640 $Y=481900
X2092 3214 3150 3141 3224 1 3205 2 AOI22S $T=542500 497400 0 0 $X=542500 $Y=497020
X2093 3219 3247 3209 2941 1 3205 2 AOI22S $T=546220 507480 1 0 $X=546220 $Y=502060
X2094 409 412 3354 410 1 411 2 AOI22S $T=564820 366360 0 0 $X=564820 $Y=365980
X2095 410 3365 3341 412 1 411 2 AOI22S $T=566060 386520 1 0 $X=566060 $Y=381100
X2096 3356 3327 3366 412 1 3360 2 AOI22S $T=566680 396600 0 0 $X=566680 $Y=396220
X2097 415 412 3359 417 1 411 2 AOI22S $T=567300 376440 1 0 $X=567300 $Y=371020
X2098 3363 3336 3362 3273 1 3346 2 AOI22S $T=567920 406680 1 0 $X=567920 $Y=401260
X2099 415 418 3344 417 1 419 2 AOI22S $T=568540 366360 0 0 $X=568540 $Y=365980
X2100 3360 417 3370 411 1 3365 2 AOI22S $T=572880 386520 1 180 $X=569160 $Y=386140
X2101 3392 3385 3399 3131 1 3316 2 AOI22S $T=574740 406680 1 180 $X=571020 $Y=406300
X2102 3346 3387 3375 3131 1 3321 2 AOI22S $T=573500 396600 1 0 $X=573500 $Y=391180
X2103 3356 3327 3404 3346 1 3273 2 AOI22S $T=574120 396600 0 0 $X=574120 $Y=396220
X2104 3392 3385 3417 3316 1 3273 2 AOI22S $T=575360 416760 1 0 $X=575360 $Y=411340
X2105 3413 3387 3412 3273 1 3356 2 AOI22S $T=579700 406680 0 180 $X=575980 $Y=401260
X2106 3363 3387 3430 3413 1 3131 2 AOI22S $T=578460 406680 0 0 $X=578460 $Y=406300
X2107 536 4002 4016 3961 1 3947 2 AOI22S $T=674560 497400 1 180 $X=670840 $Y=497020
X2108 536 4002 4018 3956 1 3983 2 AOI22S $T=675800 517560 0 180 $X=672080 $Y=512140
X2109 536 4002 4037 3927 1 3626 2 AOI22S $T=679520 497400 0 180 $X=675800 $Y=491980
X2110 536 4002 4048 3988 1 3993 2 AOI22S $T=681380 467160 0 180 $X=677660 $Y=461740
X2111 536 4002 4057 4062 1 3954 2 AOI22S $T=680760 457080 0 0 $X=680760 $Y=456700
X2112 4123 552 4112 4004 1 3801 2 AOI22S $T=693780 497400 0 180 $X=690060 $Y=491980
X2113 4097 4106 4101 4098 1 3675 2 AOI22S $T=690060 507480 0 0 $X=690060 $Y=507100
X2114 4097 4106 4088 4109 1 4046 2 AOI22S $T=690060 517560 0 0 $X=690060 $Y=517180
X2115 556 552 4124 4054 1 3707 2 AOI22S $T=696260 537720 0 180 $X=692540 $Y=532300
X2116 557 555 4122 3825 1 4013 2 AOI22S $T=696880 487320 0 180 $X=693160 $Y=481900
X2117 4123 552 4140 4039 1 4064 2 AOI22S $T=698120 497400 0 180 $X=694400 $Y=491980
X2118 4097 4131 4116 3990 1 3999 2 AOI22S $T=698740 447000 1 180 $X=695020 $Y=446620
X2119 4161 4138 4139 3928 1 4052 2 AOI22S $T=700600 426840 0 180 $X=696880 $Y=421420
X2120 4159 4152 4154 4129 1 4107 2 AOI22S $T=701840 406680 0 180 $X=698120 $Y=401260
X2121 557 555 4148 4096 1 4144 2 AOI22S $T=698120 477240 1 0 $X=698120 $Y=471820
X2122 4159 4152 4170 4095 1 4133 2 AOI22S $T=702460 416760 1 180 $X=698740 $Y=416380
X2123 4097 4106 4151 3695 1 3811 2 AOI22S $T=699360 507480 0 0 $X=699360 $Y=507100
X2124 557 555 4155 4150 1 4137 2 AOI22S $T=699980 467160 0 0 $X=699980 $Y=466780
X2125 4161 4138 4135 4160 1 4104 2 AOI22S $T=704320 436920 1 180 $X=700600 $Y=436540
X2126 4159 4152 4182 4176 1 4020 2 AOI22S $T=706180 416760 0 0 $X=706180 $Y=416380
X2127 4097 569 4165 571 1 491 2 AOI22S $T=706180 537720 1 0 $X=706180 $Y=532300
X2128 4206 575 4199 4143 1 4060 2 AOI22S $T=711760 386520 1 180 $X=708040 $Y=386140
X2129 4206 575 4211 4191 1 4079 2 AOI22S $T=714240 396600 0 180 $X=710520 $Y=391180
X2130 4206 4214 4195 581 1 4113 2 AOI22S $T=712380 386520 1 0 $X=712380 $Y=381100
X2131 4123 4216 4203 4209 1 3841 2 AOI22S $T=713000 497400 0 0 $X=713000 $Y=497020
X2132 4242 555 4208 4212 1 3765 2 AOI22S $T=717960 477240 0 180 $X=714240 $Y=471820
X2133 4206 4214 4251 4224 1 4221 2 AOI22S $T=722920 386520 1 180 $X=719200 $Y=386140
X2134 4161 4131 4253 4177 1 4072 2 AOI22S $T=723540 436920 0 180 $X=719820 $Y=431500
X2135 4123 4216 4254 4235 1 4217 2 AOI22S $T=723540 497400 0 180 $X=719820 $Y=491980
X2136 4159 4152 4264 4222 1 4227 2 AOI22S $T=725400 406680 0 180 $X=721680 $Y=401260
X2137 4242 4271 4265 4260 1 4280 2 AOI22S $T=724160 467160 0 0 $X=724160 $Y=466780
X2138 574 4106 4262 584 1 586 2 AOI22S $T=724780 527640 0 0 $X=724780 $Y=527260
X2139 4288 4281 4289 3952 1 3804 2 AOI22S $T=729120 447000 0 180 $X=725400 $Y=441580
X2140 4206 4214 4313 593 1 4294 2 AOI22S $T=734700 386520 1 180 $X=730980 $Y=386140
X2141 574 4106 4301 4293 1 587 2 AOI22S $T=730980 527640 0 0 $X=730980 $Y=527260
X2142 4242 4271 4295 4326 1 4247 2 AOI22S $T=733460 477240 1 0 $X=733460 $Y=471820
X2143 4159 4152 4310 4021 1 600 2 AOI22S $T=734700 406680 1 0 $X=734700 $Y=401260
X2144 4161 4131 4317 4287 1 4229 2 AOI22S $T=738420 436920 0 180 $X=734700 $Y=431500
X2145 4288 4281 4291 4243 1 4312 2 AOI22S $T=734700 447000 1 0 $X=734700 $Y=441580
X2146 4316 4306 4299 3742 1 4329 2 AOI22S $T=735940 497400 0 0 $X=735940 $Y=497020
X2147 4206 4214 4344 4302 1 603 2 AOI22S $T=741520 386520 0 180 $X=737800 $Y=381100
X2148 4161 4131 4384 4364 1 4352 2 AOI22S $T=748340 436920 0 180 $X=744620 $Y=431500
X2149 4288 4281 4394 4395 1 4391 2 AOI22S $T=753920 447000 0 180 $X=750200 $Y=441580
X2150 595 626 4406 625 1 4270 2 AOI22S $T=755160 537720 0 180 $X=751440 $Y=532300
X2151 4443 4433 4448 4369 1 601 2 AOI22S $T=761980 406680 1 180 $X=758260 $Y=406300
X2152 4456 4450 4453 4403 1 4373 2 AOI22S $T=765080 396600 0 180 $X=761360 $Y=391180
X2153 4441 4216 4466 4460 1 3667 2 AOI22S $T=767560 487320 1 180 $X=763840 $Y=486940
X2154 4441 4216 4472 4473 1 3739 2 AOI22S $T=766940 507480 1 0 $X=766940 $Y=502060
X2155 4242 4271 4503 4447 1 3970 2 AOI22S $T=771900 477240 0 180 $X=768180 $Y=471820
X2156 4443 4433 4485 4489 1 4499 2 AOI22S $T=769420 406680 0 0 $X=769420 $Y=406300
X2157 4443 4433 4511 4484 1 4367 2 AOI22S $T=775000 376440 1 180 $X=771280 $Y=376060
X2158 4456 4433 4497 4476 1 4519 2 AOI22S $T=771280 396600 0 0 $X=771280 $Y=396220
X2159 4462 4475 4514 4505 1 3893 2 AOI22S $T=775000 517560 0 180 $X=771280 $Y=512140
X2160 642 575 4501 631 1 647 2 AOI22S $T=771900 366360 0 0 $X=771900 $Y=365980
X2161 4462 4475 4515 3641 1 648 2 AOI22S $T=773760 517560 0 0 $X=773760 $Y=517180
X2162 4288 4281 4498 4440 1 4502 2 AOI22S $T=778100 436920 1 180 $X=774380 $Y=436540
X2163 4410 4412 4486 4506 1 4314 2 AOI22S $T=775000 416760 1 0 $X=775000 $Y=411340
X2164 4410 4412 4573 4583 1 4568 2 AOI22S $T=790500 406680 0 0 $X=790500 $Y=406300
X2165 4586 4581 4584 4579 1 4571 2 AOI22S $T=794220 477240 0 180 $X=790500 $Y=471820
X2166 618 665 4593 4602 1 4569 2 AOI22S $T=794840 376440 1 0 $X=794840 $Y=371020
X2167 618 665 4606 669 1 4601 2 AOI22S $T=797320 376440 0 0 $X=797320 $Y=376060
X2168 4578 4530 4607 4580 1 4592 2 AOI22S $T=803520 436920 0 180 $X=799800 $Y=431500
X2169 4410 4412 4632 673 1 4637 2 AOI22S $T=801660 406680 0 0 $X=801660 $Y=406300
X2170 4578 4530 4633 4644 1 676 2 AOI22S $T=802280 436920 0 0 $X=802280 $Y=436540
X2171 4586 4581 4651 4620 1 4640 2 AOI22S $T=806620 477240 0 180 $X=802900 $Y=471820
X2172 4635 4614 4636 677 1 4653 2 AOI22S $T=802900 507480 0 0 $X=802900 $Y=507100
X2173 4586 4581 4650 4656 1 4663 2 AOI22S $T=804760 467160 0 0 $X=804760 $Y=466780
X2174 4578 4530 4648 4659 1 4672 2 AOI22S $T=805380 436920 1 0 $X=805380 $Y=431500
X2175 4586 4581 4660 681 1 4673 2 AOI22S $T=806620 477240 1 0 $X=806620 $Y=471820
X2176 4667 655 4652 4012 1 685 2 AOI22S $T=807860 527640 0 0 $X=807860 $Y=527260
X2177 710 708 709 703 1 471 2 AOI22S $T=835140 537720 0 180 $X=831420 $Y=532300
X2178 4793 4778 4785 4772 1 4750 2 AOI22S $T=837620 396600 1 180 $X=833900 $Y=396220
X2179 4793 4778 4794 713 1 4691 2 AOI22S $T=838860 386520 1 180 $X=835140 $Y=386140
X2180 4793 4778 4796 716 1 715 2 AOI22S $T=839480 366360 1 180 $X=835760 $Y=365980
X2181 4793 4778 4809 4770 1 4730 2 AOI22S $T=839480 376440 1 180 $X=835760 $Y=376060
X2182 4797 4790 4815 4758 1 707 2 AOI22S $T=841340 467160 0 180 $X=837620 $Y=461740
X2183 725 708 4806 4738 1 4729 2 AOI22S $T=841340 507480 0 180 $X=837620 $Y=502060
X2184 4793 4778 727 690 1 4735 2 AOI22S $T=843200 366360 1 180 $X=839480 $Y=365980
X2185 4797 4778 4814 4784 1 4808 2 AOI22S $T=843820 406680 0 180 $X=840100 $Y=401260
X2186 4797 4790 4825 714 1 706 2 AOI22S $T=843820 426840 1 180 $X=840100 $Y=426460
X2187 4797 4790 4818 4766 1 4816 2 AOI22S $T=842580 436920 0 0 $X=842580 $Y=436540
X2188 735 736 4827 4769 1 741 2 AOI22S $T=845680 527640 0 0 $X=845680 $Y=527260
X2189 750 744 4859 726 1 4835 2 AOI22S $T=853740 507480 0 180 $X=850020 $Y=502060
X2190 4875 4865 4869 737 1 747 2 AOI22S $T=855600 376440 0 180 $X=851880 $Y=371020
X2191 4872 4858 4862 4763 1 4800 2 AOI22S $T=856220 467160 1 180 $X=852500 $Y=466780
X2192 4872 4865 4846 4836 1 4843 2 AOI22S $T=856840 426840 1 180 $X=853120 $Y=426460
X2193 4872 4865 4899 739 1 4817 2 AOI22S $T=858700 447000 1 180 $X=854980 $Y=446620
X2194 4875 4891 4877 760 1 749 2 AOI22S $T=859940 376440 0 180 $X=856220 $Y=371020
X2195 735 736 4882 4889 1 748 2 AOI22S $T=856220 507480 0 0 $X=856220 $Y=507100
X2196 4875 4865 4930 4834 1 4881 2 AOI22S $T=864900 386520 1 180 $X=861180 $Y=386140
X2197 4894 4933 4874 4908 1 4939 2 AOI22S $T=863040 396600 1 0 $X=863040 $Y=391180
X2198 4894 4903 4867 4871 1 4900 2 AOI22S $T=868000 406680 0 180 $X=864280 $Y=401260
X2199 4894 4903 4937 4929 1 4948 2 AOI22S $T=865520 447000 0 0 $X=865520 $Y=446620
X2200 4875 4891 4957 774 1 772 2 AOI22S $T=871100 376440 0 180 $X=867380 $Y=371020
X2201 4962 4955 4911 4953 1 4949 2 AOI22S $T=871100 517560 0 180 $X=867380 $Y=512140
X2202 4894 4903 4860 771 1 4950 2 AOI22S $T=869860 436920 1 0 $X=869860 $Y=431500
X2203 4894 4903 4959 4999 1 4986 2 AOI22S $T=872960 406680 0 0 $X=872960 $Y=406300
X2204 4962 4955 4864 4978 1 4952 2 AOI22S $T=876680 477240 1 180 $X=872960 $Y=476860
X2205 785 4955 4844 4987 1 4992 2 AOI22S $T=874820 426840 1 0 $X=874820 $Y=421420
X2206 785 791 4974 4984 1 793 2 AOI22S $T=875440 386520 0 0 $X=875440 $Y=386140
X2207 4962 4955 4861 4993 1 4998 2 AOI22S $T=875440 467160 1 0 $X=875440 $Y=461740
X2208 4962 779 4994 795 1 4976 2 AOI22S $T=876680 517560 1 0 $X=876680 $Y=512140
X2209 4962 4955 4914 5001 1 5003 2 AOI22S $T=877300 447000 0 0 $X=877300 $Y=446620
X2210 5008 4823 5010 4995 1 5030 2 AOI22S $T=879780 507480 1 0 $X=879780 $Y=502060
X2211 5008 5084 5088 5080 1 5078 2 AOI22S $T=897760 487320 1 180 $X=894040 $Y=486940
X2212 5089 4983 5040 5097 1 5099 2 AOI22S $T=896520 517560 1 0 $X=896520 $Y=512140
X2213 5091 4933 4981 5093 1 5111 2 AOI22S $T=899620 396600 1 0 $X=899620 $Y=391180
X2214 5091 4933 5101 5112 1 812 2 AOI22S $T=900240 396600 0 0 $X=900240 $Y=396220
X2215 5008 5084 5147 5128 1 5102 2 AOI22S $T=907060 467160 1 180 $X=903340 $Y=466780
X2216 5143 5135 5137 5113 1 5087 2 AOI22S $T=907680 426840 1 180 $X=903960 $Y=426460
X2217 5089 4983 5132 5085 1 5141 2 AOI22S $T=904580 517560 1 0 $X=904580 $Y=512140
X2218 5153 4891 5116 824 1 5142 2 AOI22S $T=910160 376440 0 180 $X=906440 $Y=371020
X2219 5163 5084 5164 814 1 5171 2 AOI22S $T=910160 457080 0 0 $X=910160 $Y=456700
X2220 5143 5084 5181 5123 1 816 2 AOI22S $T=915120 447000 1 180 $X=911400 $Y=446620
X2221 5089 4983 5195 5177 1 834 2 AOI22S $T=918220 497400 0 180 $X=914500 $Y=491980
X2222 5143 5135 5213 5108 1 5173 2 AOI22S $T=919460 436920 1 180 $X=915740 $Y=436540
X2223 757 4933 5196 5199 1 5211 2 AOI22S $T=918220 396600 0 0 $X=918220 $Y=396220
X2224 5154 5226 5246 5234 1 5186 2 AOI22S $T=926280 436920 0 180 $X=922560 $Y=431500
X2225 5143 5135 5256 5230 1 841 2 AOI22S $T=929380 416760 0 180 $X=925660 $Y=411340
X2226 5089 5226 5247 5237 1 5139 2 AOI22S $T=926900 497400 1 0 $X=926900 $Y=491980
X2227 857 5263 5051 5244 1 5257 2 AOI22S $T=932480 527640 0 180 $X=928760 $Y=522220
X2228 5153 5242 5258 854 1 861 2 AOI22S $T=929380 376440 1 0 $X=929380 $Y=371020
X2229 5143 5135 5271 5198 1 826 2 AOI22S $T=933100 386520 0 180 $X=929380 $Y=381100
X2230 5154 5226 5269 853 1 5260 2 AOI22S $T=933100 447000 0 180 $X=929380 $Y=441580
X2231 5154 5226 5275 856 1 5267 2 AOI22S $T=934340 457080 0 180 $X=930620 $Y=451660
X2232 5153 5242 5297 867 1 865 2 AOI22S $T=938060 376440 0 180 $X=934340 $Y=371020
X2233 5286 5135 5303 5264 1 868 2 AOI22S $T=938680 386520 1 180 $X=934960 $Y=386140
X2234 5154 5226 5284 5274 1 858 2 AOI22S $T=934960 457080 1 0 $X=934960 $Y=451660
X2235 5283 5289 5204 863 1 5295 2 AOI22S $T=935580 487320 0 0 $X=935580 $Y=486940
X2236 873 871 5233 5227 1 5296 2 AOI22S $T=940540 507480 0 180 $X=936820 $Y=502060
X2237 857 5289 5145 872 1 5305 2 AOI22S $T=936820 517560 0 0 $X=936820 $Y=517180
X2238 5286 5135 5298 5302 1 869 2 AOI22S $T=937440 386520 1 0 $X=937440 $Y=381100
X2239 5153 5242 5301 870 1 876 2 AOI22S $T=938680 376440 1 0 $X=938680 $Y=371020
X2240 5272 5309 5262 5311 1 5310 2 AOI22S $T=939300 416760 1 0 $X=939300 $Y=411340
X2241 873 871 5130 5339 1 887 2 AOI22S $T=944880 517560 0 0 $X=944880 $Y=517180
X2242 5272 5309 5331 886 1 890 2 AOI22S $T=945500 386520 0 0 $X=945500 $Y=386140
X2243 888 893 5316 895 1 899 2 AOI22S $T=947360 366360 0 0 $X=947360 $Y=365980
X2244 873 5344 5351 5343 1 892 2 AOI22S $T=951080 487320 1 180 $X=947360 $Y=486940
X2245 5272 5309 5352 901 1 5335 2 AOI22S $T=949840 386520 0 0 $X=949840 $Y=386140
X2246 5272 5309 5307 878 1 5359 2 AOI22S $T=949840 396600 1 0 $X=949840 $Y=391180
X2247 5354 5344 5357 891 1 898 2 AOI22S $T=953560 447000 1 180 $X=949840 $Y=446620
X2248 5354 5344 5345 5365 1 5280 2 AOI22S $T=951700 457080 0 0 $X=951700 $Y=456700
X2249 888 893 5273 902 1 903 2 AOI22S $T=952320 366360 0 0 $X=952320 $Y=365980
X2250 5283 5289 5341 905 1 5377 2 AOI22S $T=953560 497400 1 0 $X=953560 $Y=491980
X2251 5354 5344 5372 5361 1 910 2 AOI22S $T=954180 447000 0 0 $X=954180 $Y=446620
X2252 5283 5289 5251 5374 1 5340 2 AOI22S $T=954180 507480 0 0 $X=954180 $Y=507100
X2253 5283 5388 5375 5389 1 5392 2 AOI22S $T=957280 477240 1 0 $X=957280 $Y=471820
X2254 5283 5388 5349 5387 1 5401 2 AOI22S $T=959140 447000 1 0 $X=959140 $Y=441580
X2255 5283 5388 5333 5395 1 923 2 AOI22S $T=962240 457080 1 0 $X=962240 $Y=451660
X2256 5472 5462 5464 5448 1 5436 2 AOI22S $T=980840 416760 1 180 $X=977120 $Y=416380
X2257 5472 5462 5463 945 1 5430 2 AOI22S $T=982080 426840 0 180 $X=978360 $Y=421420
X2258 5481 5477 5452 927 1 947 2 AOI22S $T=983320 396600 1 180 $X=979600 $Y=396220
X2259 5481 957 5490 5441 1 5471 2 AOI22S $T=985800 497400 1 180 $X=982080 $Y=497020
X2260 5481 5477 5484 938 1 5496 2 AOI22S $T=983320 396600 0 0 $X=983320 $Y=396220
X2261 5472 5462 5499 5480 1 5488 2 AOI22S $T=987660 416760 1 180 $X=983940 $Y=416380
X2262 5512 962 5503 5493 1 5434 2 AOI22S $T=987660 457080 1 180 $X=983940 $Y=456700
X2263 5472 5462 5478 5525 1 5491 2 AOI22S $T=984560 426840 1 0 $X=984560 $Y=421420
X2264 5481 957 5498 5446 1 5528 2 AOI22S $T=985180 507480 1 0 $X=985180 $Y=502060
X2265 5481 5477 5451 968 1 972 2 AOI22S $T=987040 396600 0 0 $X=987040 $Y=396220
X2266 5495 5516 5501 974 1 5437 2 AOI22S $T=992620 477240 0 180 $X=988900 $Y=471820
X2267 5512 978 979 935 1 977 2 AOI22S $T=993860 527640 1 180 $X=990140 $Y=527260
X2268 5517 957 5543 5532 1 5552 2 AOI22S $T=995100 507480 0 0 $X=995100 $Y=507100
X2269 5495 5516 5548 5551 1 5541 2 AOI22S $T=995720 487320 1 0 $X=995720 $Y=481900
X2270 5512 978 5558 940 1 987 2 AOI22S $T=997580 527640 0 0 $X=997580 $Y=527260
X2271 5586 5567 5504 5523 1 5524 2 AOI22S $T=1001920 467160 0 180 $X=998200 $Y=461740
X2272 5517 957 5566 988 1 990 2 AOI22S $T=998820 537720 1 0 $X=998820 $Y=532300
X2273 5586 5567 5581 5610 1 5602 2 AOI22S $T=1004400 467160 1 0 $X=1004400 $Y=461740
X2274 1003 1001 5585 5606 1 997 2 AOI22S $T=1008740 376440 0 180 $X=1005020 $Y=371020
X2275 5573 5613 5582 5618 1 5633 2 AOI22S $T=1005640 416760 1 0 $X=1005640 $Y=411340
X2276 5495 5516 5595 5634 1 5564 2 AOI22S $T=1008120 426840 0 0 $X=1008120 $Y=426460
X2277 5495 5516 5625 5639 1 1008 2 AOI22S $T=1008740 487320 1 0 $X=1008740 $Y=481900
X2278 5517 5599 5593 1006 1 5609 2 AOI22S $T=1008740 507480 0 0 $X=1008740 $Y=507100
X2279 1007 1009 5605 1013 1 5624 2 AOI22S $T=1010600 527640 0 0 $X=1010600 $Y=527260
X2280 5662 5641 5520 5663 1 1019 2 AOI22S $T=1017420 487320 0 0 $X=1017420 $Y=486940
X2281 1003 1030 5688 5682 1 5660 2 AOI22S $T=1024240 406680 1 0 $X=1024240 $Y=401260
X2282 5670 1029 5590 5638 1 5706 2 AOI22S $T=1024240 527640 0 0 $X=1024240 $Y=527260
X2283 5670 1029 5693 5714 1 5702 2 AOI22S $T=1025480 487320 1 0 $X=1025480 $Y=481900
X2284 5517 5599 5704 1034 1 1033 2 AOI22S $T=1029820 507480 1 180 $X=1026100 $Y=507100
X2285 5662 5641 5710 5694 1 1041 2 AOI22S $T=1032300 497400 0 0 $X=1032300 $Y=497020
X2286 1047 5728 5730 1043 1 5729 2 AOI22S $T=1036640 447000 0 180 $X=1032920 $Y=441580
X2287 5670 5567 5720 5698 1 5735 2 AOI22S $T=1034160 467160 0 0 $X=1034160 $Y=466780
X2288 5662 5680 5725 5703 1 5747 2 AOI22S $T=1035400 426840 0 0 $X=1035400 $Y=426460
X2289 1059 5728 5715 1053 1 1052 2 AOI22S $T=1044700 366360 1 180 $X=1040980 $Y=365980
X2290 1007 5641 5778 5785 1 5793 2 AOI22S $T=1044700 517560 1 0 $X=1044700 $Y=512140
X2291 5749 5599 5792 5797 1 5736 2 AOI22S $T=1047800 497400 0 0 $X=1047800 $Y=497020
X2292 5804 5567 5805 5813 1 5791 2 AOI22S $T=1049040 477240 1 0 $X=1049040 $Y=471820
X2293 1059 5728 5824 1070 1 1072 2 AOI22S $T=1058340 376440 0 180 $X=1054620 $Y=371020
X2294 5670 5567 5827 1074 1 1075 2 AOI22S $T=1054620 467160 0 0 $X=1054620 $Y=466780
X2295 5754 5613 5838 5828 1 5801 2 AOI22S $T=1057100 406680 1 0 $X=1057100 $Y=401260
X2296 5804 5816 5891 1071 1 5752 2 AOI22S $T=1069500 477240 1 180 $X=1065780 $Y=476860
X2297 5749 5829 5897 5868 1 5833 2 AOI22S $T=1070120 497400 0 180 $X=1066400 $Y=491980
X2298 5709 5787 5893 5899 1 5890 2 AOI22S $T=1067640 447000 0 0 $X=1067640 $Y=446620
X2299 5754 5896 5925 5870 1 5874 2 AOI22S $T=1076940 406680 0 180 $X=1073220 $Y=401260
X2300 5754 5896 5943 5941 1 5920 2 AOI22S $T=1081900 396600 0 180 $X=1078180 $Y=391180
X2301 1059 1082 5940 1094 1 5948 2 AOI22S $T=1078800 376440 1 0 $X=1078800 $Y=371020
X2302 1102 5966 5954 5846 1 5909 2 AOI22S $T=1086860 517560 1 180 $X=1083140 $Y=517180
X2303 5709 5973 5964 5937 1 5968 2 AOI22S $T=1088100 457080 0 180 $X=1084380 $Y=451660
X2304 5804 5816 5962 5956 1 5928 2 AOI22S $T=1084380 467160 0 0 $X=1084380 $Y=466780
X2305 1102 5966 5971 5983 1 5960 2 AOI22S $T=1090580 517560 1 180 $X=1086860 $Y=517180
X2306 5754 5896 5984 5986 1 5995 2 AOI22S $T=1088100 396600 1 0 $X=1088100 $Y=391180
X2307 5754 5896 5981 5991 1 5997 2 AOI22S $T=1088100 406680 1 0 $X=1088100 $Y=401260
X2308 5709 5973 5944 5972 1 5992 2 AOI22S $T=1088720 447000 0 0 $X=1088720 $Y=446620
X2309 5749 5829 6025 6018 1 6016 2 AOI22S $T=1098020 497400 0 180 $X=1094300 $Y=491980
X2310 6005 5816 6039 6021 1 6030 2 AOI22S $T=1100500 477240 1 180 $X=1096780 $Y=476860
X2311 6042 5973 6050 6012 1 6038 2 AOI22S $T=1101120 447000 0 0 $X=1101120 $Y=446620
X2312 5760 6067 6000 6069 1 1119 2 AOI22S $T=1104840 406680 0 0 $X=1104840 $Y=406300
X2313 1118 1087 5961 1120 1 6059 2 AOI22S $T=1106080 366360 0 0 $X=1106080 $Y=365980
X2314 6005 5816 6066 6082 1 6079 2 AOI22S $T=1106080 477240 0 0 $X=1106080 $Y=476860
X2315 6068 5829 6065 6076 1 6064 2 AOI22S $T=1106080 497400 0 0 $X=1106080 $Y=497020
X2316 5760 6067 5963 6078 1 6095 2 AOI22S $T=1106700 416760 0 0 $X=1106700 $Y=416380
X2317 5760 6067 5976 6046 1 6108 2 AOI22S $T=1107320 406680 1 0 $X=1107320 $Y=401260
X2318 6042 5973 6053 6102 1 6105 2 AOI22S $T=1109800 447000 0 0 $X=1109800 $Y=446620
X2319 1102 5966 6077 6109 1 6056 2 AOI22S $T=1111040 527640 1 0 $X=1111040 $Y=522220
X2320 4254 4262 4272 4265 2 1 4285 AN4S $T=723540 497400 1 0 $X=723540 $Y=491980
X2321 4320 4301 4299 4295 2 1 4290 AN4S $T=734080 497400 0 180 $X=729120 $Y=491980
X2322 4383 4384 4394 4344 2 1 4409 AN4S $T=749580 436920 1 0 $X=749580 $Y=431500
X2323 4448 4457 4461 4467 2 1 4477 AN4S $T=763840 406680 0 0 $X=763840 $Y=406300
X2324 4485 4486 4498 4501 2 1 4516 AN4S $T=770040 416760 1 0 $X=770040 $Y=411340
X2325 4449 644 4512 4503 2 1 4523 AN4S $T=771900 487320 0 0 $X=771900 $Y=486940
X2326 4406 4521 4525 4528 2 1 4546 AN4S $T=775000 507480 0 0 $X=775000 $Y=507100
X2327 4453 4573 4577 661 2 1 4590 AN4S $T=789260 396600 1 0 $X=789260 $Y=391180
X2328 4472 4562 4603 4584 2 1 4616 AN4S $T=794840 507480 1 0 $X=794840 $Y=502060
X2329 4520 4599 4607 4606 2 1 4621 AN4S $T=795460 396600 1 0 $X=795460 $Y=391180
X2330 4497 4622 4633 672 2 1 4649 AN4S $T=800420 396600 0 0 $X=800420 $Y=396220
X2331 4466 4652 4657 4650 2 1 4674 AN4S $T=804760 487320 1 0 $X=804760 $Y=481900
X2332 4515 679 4636 4651 2 1 4683 AN4S $T=806000 517560 0 0 $X=806000 $Y=517180
X2333 4514 4685 4679 4660 2 1 4705 AN4S $T=812200 517560 0 0 $X=812200 $Y=517180
X2334 4860 4825 4846 4844 2 1 4710 AN4S $T=853120 426840 1 180 $X=848160 $Y=426460
X2335 4827 709 4852 4857 2 1 752 AN4S $T=849400 527640 0 0 $X=849400 $Y=527260
X2336 4887 4815 4862 4861 2 1 4839 AN4S $T=855600 467160 0 180 $X=850640 $Y=461740
X2337 4880 4795 4866 4864 2 1 4853 AN4S $T=856220 477240 1 180 $X=851260 $Y=476860
X2338 4867 4785 4877 755 2 1 4901 AN4S $T=853740 396600 0 0 $X=853740 $Y=396220
X2339 4874 4809 4869 761 2 1 4902 AN4S $T=855600 376440 0 0 $X=855600 $Y=376060
X2340 4882 4806 4859 4911 2 1 4942 AN4S $T=858080 507480 1 0 $X=858080 $Y=502060
X2341 4937 4818 4899 4914 2 1 4791 AN4S $T=864900 447000 1 180 $X=859940 $Y=446620
X2342 4959 4794 4930 4974 2 1 4985 AN4S $T=870480 386520 0 0 $X=870480 $Y=386140
X2343 4981 4796 4957 794 2 1 5012 AN4S $T=876060 376440 0 0 $X=876060 $Y=376060
X2344 5015 4814 5016 804 2 1 5032 AN4S $T=882260 396600 0 0 $X=882260 $Y=396220
X2345 5051 5010 5040 4994 2 1 5025 AN4S $T=889700 517560 0 180 $X=884740 $Y=512140
X2346 5101 727 5116 817 2 1 5100 AN4S $T=900860 376440 0 0 $X=900860 $Y=376060
X2347 5145 5070 5132 5130 2 1 5121 AN4S $T=907680 517560 1 180 $X=902720 $Y=517180
X2348 5204 5152 5195 5193 2 1 5161 AN4S $T=919460 487320 1 180 $X=914500 $Y=486940
X2349 5196 5137 5202 839 2 1 5221 AN4S $T=916980 396600 1 0 $X=916980 $Y=391180
X2350 5251 5088 5231 5233 2 1 5188 AN4S $T=926900 507480 0 180 $X=921940 $Y=502060
X2351 5262 5256 5246 5273 2 1 5291 AN4S $T=930620 416760 1 0 $X=930620 $Y=411340
X2352 5307 5303 5258 5316 2 1 5326 AN4S $T=939920 386520 0 0 $X=939920 $Y=386140
X2353 5333 5181 5284 5345 2 1 5353 AN4S $T=946120 457080 1 0 $X=946120 $Y=451660
X2354 5331 5271 5297 897 2 1 5358 AN4S $T=947980 386520 1 0 $X=947980 $Y=381100
X2355 5341 5147 5247 5351 2 1 5362 AN4S $T=947980 497400 1 0 $X=947980 $Y=491980
X2356 5349 5213 5269 5357 2 1 5367 AN4S $T=949840 447000 1 0 $X=949840 $Y=441580
X2357 5352 5298 5301 906 2 1 5382 AN4S $T=952940 386520 1 0 $X=952940 $Y=381100
X2358 5375 5164 5275 5372 2 1 5399 AN4S $T=956040 457080 1 0 $X=956040 $Y=451660
X2359 5566 5605 5558 5590 2 1 994 AN4S $T=1006880 527640 1 180 $X=1001920 $Y=527260
X2360 5704 5712 5693 5710 2 1 4783 AN4S $T=1032300 497400 0 180 $X=1027340 $Y=491980
X2361 5726 5732 5688 5725 2 1 4707 AN4S $T=1035400 406680 0 180 $X=1030440 $Y=401260
X2362 5792 5778 5784 5805 2 1 4854 AN4S $T=1046560 487320 1 0 $X=1046560 $Y=481900
X2363 5838 5830 5824 1069 2 1 5009 AN4S $T=1056480 406680 0 180 $X=1051520 $Y=401260
X2364 5897 5877 5893 5891 2 1 4868 AN4S $T=1070740 487320 0 180 $X=1065780 $Y=481900
X2365 5933 5954 5944 5942 2 1 5115 AN4S $T=1083140 497400 0 180 $X=1078180 $Y=491980
X2366 5925 5963 1099 1098 2 1 5029 AN4S $T=1085620 406680 1 180 $X=1080660 $Y=406300
X2367 5981 5970 1101 5961 2 1 5005 AN4S $T=1086860 406680 0 180 $X=1081900 $Y=401260
X2368 5982 5971 5964 5962 2 1 5165 AN4S $T=1086860 487320 1 180 $X=1081900 $Y=486940
X2369 5984 6000 1105 5989 2 1 5002 AN4S $T=1092440 386520 0 180 $X=1087480 $Y=381100
X2370 6065 6058 6053 6052 2 1 4936 AN4S $T=1105460 497400 1 180 $X=1100500 $Y=497020
X2371 1205 2 1 11 BUF1 $T=220720 366360 0 0 $X=220720 $Y=365980
X2372 8 2 1 3 BUF1 $T=223200 416760 1 180 $X=220720 $Y=416380
X2373 1234 2 1 1219 BUF1 $T=226300 507480 0 180 $X=223820 $Y=502060
X2374 1243 2 1 15 BUF1 $T=228160 497400 1 180 $X=225680 $Y=497020
X2375 1250 2 1 17 BUF1 $T=230020 467160 1 180 $X=227540 $Y=466780
X2376 25 2 1 1217 BUF1 $T=228160 497400 0 0 $X=228160 $Y=497020
X2377 1296 2 1 1278 BUF1 $T=238080 507480 1 0 $X=238080 $Y=502060
X2378 1234 2 1 1319 BUF1 $T=239940 517560 1 0 $X=239940 $Y=512140
X2379 38 2 1 24 BUF1 $T=243040 507480 0 180 $X=240560 $Y=502060
X2380 45 2 1 1305 BUF1 $T=247380 527640 1 0 $X=247380 $Y=522220
X2381 1305 2 1 1359 BUF1 $T=249240 507480 0 0 $X=249240 $Y=507100
X2382 1319 2 1 51 BUF1 $T=249240 527640 0 0 $X=249240 $Y=527260
X2383 50 2 1 32 BUF1 $T=252960 497400 1 180 $X=250480 $Y=497020
X2384 1835 2 1 1674 BUF1 $T=326740 507480 0 180 $X=324260 $Y=502060
X2385 135 2 1 1853 BUF1 $T=346580 447000 0 0 $X=346580 $Y=446620
X2386 2106 2 1 2098 BUF1 $T=373240 467160 0 0 $X=373240 $Y=466780
X2387 2187 2 1 2106 BUF1 $T=388120 457080 0 180 $X=385640 $Y=451660
X2388 2182 2 1 2245 BUF1 $T=393700 457080 0 0 $X=393700 $Y=456700
X2389 2032 2 1 2222 BUF1 $T=395560 477240 0 0 $X=395560 $Y=476860
X2390 188 2 1 2032 BUF1 $T=396180 487320 0 0 $X=396180 $Y=486940
X2391 2222 2 1 2119 BUF1 $T=398040 436920 0 0 $X=398040 $Y=436540
X2392 195 2 1 2145 BUF1 $T=401140 386520 0 180 $X=398660 $Y=381100
X2393 2280 2 1 1837 BUF1 $T=403000 487320 1 180 $X=400520 $Y=486940
X2394 2260 2 1 186 BUF1 $T=401140 426840 0 0 $X=401140 $Y=426460
X2395 198 2 1 2251 BUF1 $T=401760 366360 0 0 $X=401760 $Y=365980
X2396 182 2 1 2128 BUF1 $T=403620 426840 0 0 $X=403620 $Y=426460
X2397 2245 2 1 196 BUF1 $T=406100 447000 0 180 $X=403620 $Y=441580
X2398 2194 2 1 2267 BUF1 $T=407960 467160 1 180 $X=405480 $Y=466780
X2399 2184 2 1 2292 BUF1 $T=407960 487320 1 180 $X=405480 $Y=486940
X2400 2267 2 1 205 BUF1 $T=406720 376440 0 0 $X=406720 $Y=376060
X2401 2317 2 1 2298 BUF1 $T=407340 447000 1 0 $X=407340 $Y=441580
X2402 2292 2 1 2181 BUF1 $T=411680 426840 1 180 $X=409200 $Y=426460
X2403 2282 2 1 2187 BUF1 $T=412920 447000 0 180 $X=410440 $Y=441580
X2404 206 2 1 2190 BUF1 $T=414780 406680 0 180 $X=412300 $Y=401260
X2405 2414 2 1 218 BUF1 $T=426560 416760 1 180 $X=424080 $Y=416380
X2406 226 2 1 220 BUF1 $T=429040 376440 0 180 $X=426560 $Y=371020
X2407 2415 2 1 224 BUF1 $T=426560 396600 0 0 $X=426560 $Y=396220
X2408 241 2 1 244 BUF1 $T=437720 366360 0 0 $X=437720 $Y=365980
X2409 2519 2 1 2518 BUF1 $T=442680 447000 1 0 $X=442680 $Y=441580
X2410 2529 2 1 241 BUF1 $T=445780 376440 1 180 $X=443300 $Y=376060
X2411 2526 2 1 254 BUF1 $T=443920 366360 0 0 $X=443920 $Y=365980
X2412 2537 2 1 2526 BUF1 $T=447020 416760 1 0 $X=447020 $Y=411340
X2413 2590 2 1 263 BUF1 $T=456940 416760 1 180 $X=454460 $Y=416380
X2414 263 2 1 266 BUF1 $T=455080 396600 0 0 $X=455080 $Y=396220
X2415 313 2 1 305 BUF1 $T=487940 477240 0 0 $X=487940 $Y=476860
X2416 2585 2 1 321 BUF1 $T=492280 487320 0 0 $X=492280 $Y=486940
X2417 2830 2 1 2585 BUF1 $T=494760 467160 1 0 $X=494760 $Y=461740
X2418 2989 2 1 2906 BUF1 $T=520180 436920 1 0 $X=520180 $Y=431500
X2419 337 2 1 3154 BUF1 $T=531960 527640 1 0 $X=531960 $Y=522220
X2420 313 2 1 3223 BUF1 $T=553040 477240 0 0 $X=553040 $Y=476860
X2421 402 2 1 3317 BUF1 $T=554900 537720 1 0 $X=554900 $Y=532300
X2422 416 2 1 3418 BUF1 $T=574120 507480 0 0 $X=574120 $Y=507100
X2423 3159 2 1 433 BUF1 $T=578460 517560 1 180 $X=575980 $Y=517180
X2424 3428 2 1 3441 BUF1 $T=577840 416760 0 0 $X=577840 $Y=416380
X2425 3159 2 1 3338 BUF1 $T=581560 487320 1 180 $X=579080 $Y=486940
X2426 3441 2 1 440 BUF1 $T=585280 366360 0 0 $X=585280 $Y=365980
X2427 447 2 1 3244 BUF1 $T=587140 527640 0 0 $X=587140 $Y=527260
X2428 3244 2 1 3608 BUF1 $T=603880 477240 0 0 $X=603880 $Y=476860
X2429 444 2 1 3614 BUF1 $T=611940 497400 0 180 $X=609460 $Y=491980
X2430 423 2 1 3630 BUF1 $T=611320 487320 0 0 $X=611320 $Y=486940
X2431 453 2 1 3658 BUF1 $T=613180 497400 1 0 $X=613180 $Y=491980
X2432 3659 2 1 3429 BUF1 $T=613800 507480 0 0 $X=613800 $Y=507100
X2433 469 2 1 3659 BUF1 $T=615660 527640 0 0 $X=615660 $Y=527260
X2434 450 2 1 3666 BUF1 $T=616280 477240 1 0 $X=616280 $Y=471820
X2435 3775 2 1 474 BUF1 $T=633640 366360 1 180 $X=631160 $Y=365980
X2436 3775 2 1 3776 BUF1 $T=634880 376440 0 0 $X=634880 $Y=376060
X2437 3823 2 1 498 BUF1 $T=651620 386520 1 180 $X=649140 $Y=386140
X2438 3916 2 1 519 BUF1 $T=661540 376440 0 0 $X=661540 $Y=376060
X2439 519 2 1 512 BUF1 $T=664640 376440 1 0 $X=664640 $Y=371020
X2440 3984 2 1 525 BUF1 $T=670840 426840 1 0 $X=670840 $Y=421420
X2441 3917 2 1 538 BUF1 $T=673940 396600 0 0 $X=673940 $Y=396220
X2442 537 2 1 3894 BUF1 $T=674560 386520 0 0 $X=674560 $Y=386140
X2443 549 2 1 4103 BUF1 $T=691300 457080 0 0 $X=691300 $Y=456700
X2444 548 2 1 4070 BUF1 $T=699360 467160 1 180 $X=696880 $Y=466780
X2445 4097 2 1 4161 BUF1 $T=697500 436920 0 0 $X=697500 $Y=436540
X2446 4106 2 1 4131 BUF1 $T=703080 457080 0 180 $X=700600 $Y=451660
X2447 566 2 1 4179 BUF1 $T=703700 517560 1 0 $X=703700 $Y=512140
X2448 574 2 1 4097 BUF1 $T=708660 527640 0 0 $X=708660 $Y=527260
X2449 4240 2 1 4245 BUF1 $T=719200 447000 1 0 $X=719200 $Y=441580
X2450 4073 2 1 4263 BUF1 $T=721680 447000 1 0 $X=721680 $Y=441580
X2451 4255 2 1 4240 BUF1 $T=724160 457080 1 180 $X=721680 $Y=456700
X2452 589 2 1 4228 BUF1 $T=730980 527640 1 180 $X=728500 $Y=527260
X2453 4228 2 1 4315 BUF1 $T=731600 487320 0 0 $X=731600 $Y=486940
X2454 595 2 1 4123 BUF1 $T=734700 497400 1 180 $X=732220 $Y=497020
X2455 599 2 1 4351 BUF1 $T=739040 527640 1 0 $X=739040 $Y=522220
X2456 4351 2 1 4255 BUF1 $T=744620 487320 1 180 $X=742140 $Y=486940
X2457 557 2 1 618 BUF1 $T=750820 457080 1 180 $X=748340 $Y=456700
X2458 4131 2 1 4412 BUF1 $T=752680 426840 0 0 $X=752680 $Y=426460
X2459 595 2 1 4441 BUF1 $T=763840 487320 1 180 $X=761360 $Y=486940
X2460 595 2 1 4462 BUF1 $T=762600 517560 1 0 $X=762600 $Y=512140
X2461 595 2 1 4443 BUF1 $T=766940 457080 1 180 $X=764460 $Y=456700
X2462 4443 2 1 4456 BUF1 $T=770040 396600 1 180 $X=767560 $Y=396220
X2463 645 2 1 4399 BUF1 $T=775000 477240 1 0 $X=775000 $Y=471820
X2464 613 2 1 4459 BUF1 $T=777480 517560 0 0 $X=777480 $Y=517180
X2465 4316 2 1 4288 BUF1 $T=778100 436920 0 0 $X=778100 $Y=436540
X2466 651 2 1 4316 BUF1 $T=784300 497400 0 180 $X=781820 $Y=491980
X2467 652 2 1 4306 BUF1 $T=784920 507480 0 180 $X=782440 $Y=502060
X2468 4530 2 1 4281 BUF1 $T=787400 436920 1 180 $X=784920 $Y=436540
X2469 4464 2 1 4518 BUF1 $T=785540 447000 0 0 $X=785540 $Y=446620
X2470 4316 2 1 4578 BUF1 $T=789260 436920 1 0 $X=789260 $Y=431500
X2471 4271 2 1 4581 BUF1 $T=797320 467160 1 180 $X=794840 $Y=466780
X2472 652 2 1 4614 BUF1 $T=796080 497400 0 0 $X=796080 $Y=497020
X2473 670 2 1 4423 BUF1 $T=798560 527640 0 0 $X=798560 $Y=527260
X2474 4610 2 1 4631 BUF1 $T=799800 406680 1 0 $X=799800 $Y=401260
X2475 653 2 1 4667 BUF1 $T=805380 527640 0 0 $X=805380 $Y=527260
X2476 686 2 1 4555 BUF1 $T=810340 507480 1 0 $X=810340 $Y=502060
X2477 4682 2 1 4695 BUF1 $T=810960 406680 1 0 $X=810960 $Y=401260
X2478 4695 2 1 4429 BUF1 $T=815300 376440 0 180 $X=812820 $Y=371020
X2479 4631 2 1 4550 BUF1 $T=815920 386520 1 180 $X=813440 $Y=386140
X2480 4315 2 1 4732 BUF1 $T=820880 436920 1 0 $X=820880 $Y=431500
X2481 725 2 1 4797 BUF1 $T=841340 497400 1 180 $X=838860 $Y=497020
X2482 684 2 1 729 BUF1 $T=840720 386520 1 0 $X=840720 $Y=381100
X2483 708 2 1 4823 BUF1 $T=841340 507480 1 0 $X=841340 $Y=502060
X2484 4790 2 1 4778 BUF1 $T=843820 406680 1 0 $X=843820 $Y=401260
X2485 731 2 1 4737 BUF1 $T=846300 477240 0 180 $X=843820 $Y=471820
X2486 721 2 1 722 BUF1 $T=843820 537720 1 0 $X=843820 $Y=532300
X2487 708 2 1 4790 BUF1 $T=845680 507480 1 0 $X=845680 $Y=502060
X2488 744 2 1 4865 BUF1 $T=851260 497400 0 0 $X=851260 $Y=497020
X2489 4255 2 1 4917 BUF1 $T=856840 457080 0 0 $X=856840 $Y=456700
X2490 777 2 1 4757 BUF1 $T=866760 436920 1 180 $X=864280 $Y=436540
X2491 757 2 1 4894 BUF1 $T=868000 436920 0 0 $X=868000 $Y=436540
X2492 744 2 1 4983 BUF1 $T=871100 507480 1 0 $X=871100 $Y=502060
X2493 776 2 1 4962 BUF1 $T=872340 537720 1 0 $X=872340 $Y=532300
X2494 4962 2 1 785 BUF1 $T=872960 426840 0 0 $X=872960 $Y=426460
X2495 4903 2 1 4933 BUF1 $T=873580 406680 1 0 $X=873580 $Y=401260
X2496 779 2 1 4955 BUF1 $T=876680 517560 1 180 $X=874200 $Y=517180
X2497 777 2 1 4970 BUF1 $T=878540 447000 0 180 $X=876060 $Y=441580
X2498 725 2 1 5008 BUF1 $T=876060 507480 1 0 $X=876060 $Y=502060
X2499 750 2 1 4941 BUF1 $T=877920 497400 0 0 $X=877920 $Y=497020
X2500 4737 2 1 797 BUF1 $T=885980 406680 1 0 $X=885980 $Y=401260
X2501 4823 2 1 5084 BUF1 $T=897760 487320 0 0 $X=897760 $Y=486940
X2502 4941 2 1 5089 BUF1 $T=904580 497400 0 0 $X=904580 $Y=497020
X2503 5084 2 1 5135 BUF1 $T=913260 436920 0 0 $X=913260 $Y=436540
X2504 4695 2 1 827 BUF1 $T=915120 396600 0 0 $X=915120 $Y=396220
X2505 4983 2 1 5226 BUF1 $T=920700 487320 0 0 $X=920700 $Y=486940
X2506 857 2 1 5283 BUF1 $T=933100 507480 1 0 $X=933100 $Y=502060
X2507 5327 2 1 844 BUF1 $T=944880 386520 1 0 $X=944880 $Y=381100
X2508 4933 2 1 5309 BUF1 $T=944880 396600 0 0 $X=944880 $Y=396220
X2509 2465 2 1 885 BUF1 $T=945500 426840 0 0 $X=945500 $Y=426460
X2510 873 2 1 5354 BUF1 $T=954800 477240 1 180 $X=952320 $Y=476860
X2511 5378 2 1 5125 BUF1 $T=957900 467160 0 180 $X=955420 $Y=461740
X2512 5045 2 1 5410 BUF1 $T=961620 517560 0 0 $X=961620 $Y=517180
X2513 864 2 1 5413 BUF1 $T=980220 507480 0 0 $X=980220 $Y=507100
X2514 956 2 1 904 BUF1 $T=985180 447000 1 180 $X=982700 $Y=446620
X2515 5495 2 1 5472 BUF1 $T=985180 426840 0 0 $X=985180 $Y=426460
X2516 962 2 1 5519 BUF1 $T=987660 457080 0 0 $X=987660 $Y=456700
X2517 5516 2 1 5462 BUF1 $T=990760 426840 0 180 $X=988280 $Y=421420
X2518 5327 2 1 976 BUF1 $T=992000 396600 1 0 $X=992000 $Y=391180
X2519 5240 2 1 5554 BUF1 $T=995720 406680 1 0 $X=995720 $Y=401260
X2520 5378 2 1 5579 BUF1 $T=1002540 457080 0 0 $X=1002540 $Y=456700
X2521 5613 2 1 5477 BUF1 $T=1008120 406680 1 180 $X=1005640 $Y=406300
X2522 931 2 1 5601 BUF1 $T=1008120 497400 1 0 $X=1008120 $Y=491980
X2523 5641 2 1 5516 BUF1 $T=1011840 477240 1 180 $X=1009360 $Y=476860
X2524 1005 2 1 5652 BUF1 $T=1016180 497400 1 0 $X=1016180 $Y=491980
X2525 1023 2 1 5668 BUF1 $T=1024860 406680 0 0 $X=1024860 $Y=406300
X2526 5567 2 1 1030 BUF1 $T=1027960 406680 1 0 $X=1027960 $Y=401260
X2527 5517 2 1 5573 BUF1 $T=1029200 426840 0 0 $X=1029200 $Y=426460
X2528 1007 2 1 5662 BUF1 $T=1029820 497400 0 0 $X=1029820 $Y=497020
X2529 5519 2 1 5728 BUF1 $T=1030440 447000 0 0 $X=1030440 $Y=446620
X2530 1029 2 1 5567 BUF1 $T=1032300 477240 0 0 $X=1032300 $Y=476860
X2531 5512 2 1 1047 BUF1 $T=1034160 447000 0 0 $X=1034160 $Y=446620
X2532 1021 2 1 5742 BUF1 $T=1034160 517560 1 0 $X=1034160 $Y=512140
X2533 5662 2 1 5760 BUF1 $T=1035400 426840 1 0 $X=1035400 $Y=421420
X2534 5573 2 1 5754 BUF1 $T=1036020 406680 0 0 $X=1036020 $Y=406300
X2535 5517 2 1 5749 BUF1 $T=1036020 497400 0 0 $X=1036020 $Y=497020
X2536 5512 2 1 5709 BUF1 $T=1037880 447000 0 0 $X=1037880 $Y=446620
X2537 1054 2 1 5613 BUF1 $T=1043460 467160 1 180 $X=1040980 $Y=466780
X2538 1054 2 1 5599 BUF1 $T=1041600 517560 1 0 $X=1041600 $Y=512140
X2539 1047 2 1 1059 BUF1 $T=1044700 366360 0 0 $X=1044700 $Y=365980
X2540 5670 2 1 5804 BUF1 $T=1045940 477240 1 0 $X=1045940 $Y=471820
X2541 1065 2 1 1063 BUF1 $T=1048420 406680 0 0 $X=1048420 $Y=406300
X2542 1029 2 1 5816 BUF1 $T=1049660 477240 0 0 $X=1049660 $Y=476860
X2543 5599 2 1 5829 BUF1 $T=1052140 497400 0 0 $X=1052140 $Y=497020
X2544 1077 2 1 1065 BUF1 $T=1058340 537720 0 180 $X=1055860 $Y=532300
X2545 5728 2 1 1082 BUF1 $T=1058960 376440 1 0 $X=1058960 $Y=371020
X2546 1080 2 1 5847 BUF1 $T=1063920 497400 1 0 $X=1063920 $Y=491980
X2547 5847 2 1 1095 BUF1 $T=1076940 416760 0 0 $X=1076940 $Y=416380
X2548 1080 2 1 1097 BUF1 $T=1079420 537720 1 0 $X=1079420 $Y=532300
X2549 1093 2 1 5911 BUF1 $T=1083140 497400 1 0 $X=1083140 $Y=491980
X2550 5519 2 1 5973 BUF1 $T=1088100 457080 1 0 $X=1088100 $Y=451660
X2551 5804 2 1 6005 BUF1 $T=1088100 467160 0 0 $X=1088100 $Y=466780
X2552 1104 2 1 5918 BUF1 $T=1090580 457080 1 0 $X=1090580 $Y=451660
X2553 5918 2 1 6043 BUF1 $T=1101740 406680 0 0 $X=1101740 $Y=406300
X2554 6080 2 1 6074 BUF1 $T=1119720 507480 1 180 $X=1117240 $Y=507100
X2555 108 1 2 1766 BUF1CK $T=316200 467160 1 0 $X=316200 $Y=461740
X2556 1850 1 2 1836 BUF1CK $T=334800 426840 1 0 $X=334800 $Y=421420
X2557 2186 1 2 179 BUF1CK $T=393080 406680 1 180 $X=390600 $Y=406300
X2558 2409 1 2 2422 BUF1CK $T=424700 477240 1 0 $X=424700 $Y=471820
X2559 2618 1 2 2629 BUF1CK $T=459420 507480 0 0 $X=459420 $Y=507100
X2560 2666 1 2 2617 BUF1CK $T=469960 477240 0 0 $X=469960 $Y=476860
X2561 2802 1 2 2734 BUF1CK $T=497240 396600 0 0 $X=497240 $Y=396220
X2562 2883 1 2 2894 BUF1CK $T=502200 386520 1 0 $X=502200 $Y=381100
X2563 2821 1 2 2953 BUF1CK $T=510260 386520 1 0 $X=510260 $Y=381100
X2564 2833 1 2 2952 BUF1CK $T=520180 366360 0 0 $X=520180 $Y=365980
X2565 2974 1 2 3056 BUF1CK $T=520800 406680 0 0 $X=520800 $Y=406300
X2566 342 1 2 3100 BUF1CK $T=525140 366360 0 0 $X=525140 $Y=365980
X2567 3094 1 2 3102 BUF1CK $T=527000 406680 1 0 $X=527000 $Y=401260
X2568 3104 1 2 3041 BUF1CK $T=527620 467160 0 0 $X=527620 $Y=466780
X2569 3163 1 2 3174 BUF1CK $T=535060 447000 1 0 $X=535060 $Y=441580
X2570 2874 1 2 3114 BUF1CK $T=541260 386520 0 0 $X=541260 $Y=386140
X2571 3126 1 2 3177 BUF1CK $T=541260 477240 0 0 $X=541260 $Y=476860
X2572 3232 1 2 3228 BUF1CK $T=547460 517560 1 0 $X=547460 $Y=512140
X2573 3295 1 2 374 BUF1CK $T=556760 467160 1 0 $X=556760 $Y=461740
X2574 2982 1 2 3281 BUF1CK $T=556760 497400 1 0 $X=556760 $Y=491980
X2575 3310 1 2 3372 BUF1CK $T=565440 487320 1 0 $X=565440 $Y=481900
X2576 416 1 2 3310 BUF1CK $T=568540 517560 1 0 $X=568540 $Y=512140
X2577 3706 1 2 485 BUF1CK $T=634880 396600 1 0 $X=634880 $Y=391180
X2578 569 1 2 4106 BUF1CK $T=706180 527640 1 180 $X=703700 $Y=527260
X2579 4327 1 2 4328 BUF1CK $T=735320 386520 1 0 $X=735320 $Y=381100
X2580 652 1 2 4530 BUF1CK $T=783060 487320 0 180 $X=780580 $Y=481900
X2581 864 1 2 5167 BUF1CK $T=959140 426840 0 0 $X=959140 $Y=426460
X2582 5406 1 2 5405 BUF1CK $T=962240 477240 0 0 $X=962240 $Y=476860
X2583 5320 1 2 5416 BUF1CK $T=968440 436920 0 0 $X=968440 $Y=436540
X2584 5538 1 2 986 BUF1CK $T=995720 537720 1 0 $X=995720 $Y=532300
X2585 864 1 2 5588 BUF1CK $T=1000680 436920 1 0 $X=1000680 $Y=431500
X2586 1004 1 2 1005 BUF1CK $T=1007500 527640 0 0 $X=1007500 $Y=527260
X2587 5662 1 2 5495 BUF1CK $T=1018040 426840 0 0 $X=1018040 $Y=426460
X2588 5746 1 2 5737 BUF1CK $T=1037880 537720 1 0 $X=1037880 $Y=532300
X2589 1058 1 2 1067 BUF1CK $T=1058340 527640 1 180 $X=1055860 $Y=527260
X2590 5410 1 2 5969 BUF1CK $T=1093060 467160 0 0 $X=1093060 $Y=466780
X2591 5709 1 2 6042 BUF1CK $T=1098020 447000 0 0 $X=1098020 $Y=446620
X2592 5749 1 2 6068 BUF1CK $T=1104220 497400 1 0 $X=1104220 $Y=491980
X2593 1233 1241 1 2 INV2 $T=228160 487320 1 0 $X=228160 $Y=481900
X2594 1287 1293 1 2 INV2 $T=234980 507480 0 0 $X=234980 $Y=507100
X2595 2558 242 1 2 INV2 $T=458180 416760 1 0 $X=458180 $Y=411340
X2596 2672 277 1 2 INV2 $T=468100 406680 0 0 $X=468100 $Y=406300
X2597 308 2519 1 2 INV2 $T=487320 527640 0 180 $X=485460 $Y=522220
X2598 2797 309 1 2 INV2 $T=489180 376440 0 180 $X=487320 $Y=371020
X2599 349 312 1 2 INV2 $T=518320 537720 0 180 $X=516460 $Y=532300
X2600 349 3159 1 2 INV2 $T=539400 527640 1 0 $X=539400 $Y=522220
X2601 3154 3305 1 2 INV2 $T=559240 477240 0 0 $X=559240 $Y=476860
X2602 3323 403 1 2 INV2 $T=560480 537720 1 0 $X=560480 $Y=532300
X2603 2982 3329 1 2 INV2 $T=565440 497400 0 0 $X=565440 $Y=497020
X2604 3329 3368 1 2 INV2 $T=568540 497400 0 0 $X=568540 $Y=497020
X2605 406 3408 1 2 INV2 $T=574120 517560 1 0 $X=574120 $Y=512140
X2606 3394 416 1 2 INV2 $T=574120 517560 0 0 $X=574120 $Y=517180
X2607 2830 437 1 2 INV2 $T=584040 467160 0 0 $X=584040 $Y=466780
X2608 407 453 1 2 INV2 $T=592100 507480 0 0 $X=592100 $Y=507100
X2609 3126 444 1 2 INV2 $T=602640 487320 0 0 $X=602640 $Y=486940
X2610 3761 3706 1 2 INV2 $T=633020 426840 0 0 $X=633020 $Y=426460
X2611 487 3775 1 2 INV2 $T=636740 366360 1 180 $X=634880 $Y=365980
X2612 3807 492 1 2 INV2 $T=638600 436920 1 180 $X=636740 $Y=436540
X2613 3877 3823 1 2 INV2 $T=649140 436920 1 180 $X=647280 $Y=436540
X2614 3863 502 1 2 INV2 $T=647900 376440 1 0 $X=647900 $Y=371020
X2615 3859 503 1 2 INV2 $T=649140 517560 0 0 $X=649140 $Y=517180
X2616 3895 505 1 2 INV2 $T=654100 376440 0 180 $X=652240 $Y=371020
X2617 3922 3917 1 2 INV2 $T=656580 467160 0 180 $X=654720 $Y=461740
X2618 3934 3916 1 2 INV2 $T=659680 467160 0 180 $X=657820 $Y=461740
X2619 3962 3984 1 2 INV2 $T=662780 447000 1 0 $X=662780 $Y=441580
X2620 2465 591 1 2 INV2 $T=732840 426840 0 0 $X=732840 $Y=426460
X2621 5278 5289 1 2 INV2 $T=943020 527640 1 0 $X=943020 $Y=522220
X2622 5440 5327 1 2 INV2 $T=972160 457080 0 0 $X=972160 $Y=456700
X2623 964 5517 1 2 INV2 $T=987040 527640 0 0 $X=987040 $Y=527260
X2624 5669 1003 1 2 INV2 $T=1020520 406680 1 180 $X=1018660 $Y=406300
X2625 1024 5670 1 2 INV2 $T=1021760 527640 0 0 $X=1021760 $Y=527260
X2626 1076 5641 1 2 INV2 $T=1058340 527640 1 0 $X=1058340 $Y=522220
X2627 1009 1076 1 2 INV2 $T=1058960 527640 0 0 $X=1058960 $Y=527260
X2628 6019 6067 1 2 INV2 $T=1104840 416760 0 0 $X=1104840 $Y=416380
X2629 218 227 1 2 BUF2 $T=429660 416760 1 0 $X=429660 $Y=411340
X2630 3074 3111 1 2 BUF2 $T=527620 447000 1 0 $X=527620 $Y=441580
X2631 3323 2982 1 2 BUF2 $T=559860 507480 0 0 $X=559860 $Y=507100
X2632 3054 407 1 2 BUF2 $T=559860 517560 1 0 $X=559860 $Y=512140
X2633 3126 346 1 2 BUF2 $T=567300 507480 0 180 $X=564200 $Y=502060
X2634 365 405 1 2 BUF2 $T=569780 527640 0 0 $X=569780 $Y=527260
X2635 3754 489 1 2 BUF2 $T=639840 376440 0 180 $X=636740 $Y=371020
X2636 3831 497 1 2 BUF2 $T=642320 376440 0 0 $X=642320 $Y=376060
X2637 3921 3920 1 2 BUF2 $T=661540 416760 1 0 $X=661540 $Y=411340
X2638 3932 528 1 2 BUF2 $T=673320 426840 1 0 $X=673320 $Y=421420
X2639 4271 575 1 2 BUF2 $T=727880 467160 0 0 $X=727880 $Y=466780
X2640 555 4271 1 2 BUF2 $T=730360 477240 1 0 $X=730360 $Y=471820
X2641 4459 4407 1 2 BUF2 $T=764460 447000 1 0 $X=764460 $Y=441580
X2642 4242 4586 1 2 BUF2 $T=794220 477240 1 0 $X=794220 $Y=471820
X2643 4865 4891 1 2 BUF2 $T=863040 376440 1 0 $X=863040 $Y=371020
X2644 722 5045 1 2 BUF2 $T=884740 527640 1 0 $X=884740 $Y=522220
X2645 825 5320 1 2 BUF2 $T=942400 447000 1 0 $X=942400 $Y=441580
X2646 982 5512 1 2 BUF2 $T=995720 537720 0 180 $X=992620 $Y=532300
X2647 5602 5568 1 2 BUF2 $T=1005020 467160 0 0 $X=1005020 $Y=466780
X2648 1003 1028 1 2 BUF2 $T=1023620 376440 1 0 $X=1023620 $Y=371020
X2649 1093 5856 1 2 BUF2 $T=1075080 396600 1 0 $X=1075080 $Y=391180
X2650 1093 5895 1 2 BUF2 $T=1081280 457080 1 0 $X=1081280 $Y=451660
X2651 5969 1115 1 2 BUF2 $T=1101120 416760 0 0 $X=1101120 $Y=416380
X2652 146 1 1979 1982 2 150 ND3 $T=354640 376440 1 0 $X=354640 $Y=371020
X2653 2808 1 2803 2810 2 281 ND3 $T=491660 436920 1 180 $X=489180 $Y=436540
X2654 2823 1 2809 2808 2 2837 ND3 $T=494140 436920 0 0 $X=494140 $Y=436540
X2655 2763 1 2875 2879 2 2811 ND3 $T=504060 416760 0 180 $X=501580 $Y=411340
X2656 2943 1 2929 2927 2 2923 ND3 $T=510880 396600 0 180 $X=508400 $Y=391180
X2657 2960 1 2985 2762 2 2996 ND3 $T=513980 386520 0 0 $X=513980 $Y=386140
X2658 3043 1 2988 2987 2 3030 ND3 $T=518320 416760 1 0 $X=518320 $Y=411340
X2659 3068 1 3072 3062 2 3132 ND3 $T=524520 406680 0 0 $X=524520 $Y=406300
X2660 3080 1 3096 3098 2 3138 ND3 $T=526380 487320 0 0 $X=526380 $Y=486940
X2661 3118 1 3127 3129 2 2994 ND3 $T=529480 507480 1 0 $X=529480 $Y=502060
X2662 3136 1 3141 3125 2 3147 ND3 $T=531340 487320 1 0 $X=531340 $Y=481900
X2663 3146 1 3140 3171 2 3155 ND3 $T=533200 396600 0 0 $X=533200 $Y=396220
X2664 3145 1 3152 3156 2 3165 ND3 $T=533200 406680 0 0 $X=533200 $Y=406300
X2665 3172 1 3167 3021 2 3087 ND3 $T=537540 376440 0 180 $X=535060 $Y=371020
X2666 381 1 3178 2829 2 380 ND3 $T=539400 366360 1 180 $X=536920 $Y=365980
X2667 382 1 3188 2840 2 3200 ND3 $T=538780 376440 1 0 $X=538780 $Y=371020
X2668 3183 1 3184 3197 2 3196 ND3 $T=538780 487320 0 0 $X=538780 $Y=486940
X2669 3189 1 3206 3210 2 3194 ND3 $T=540640 416760 0 0 $X=540640 $Y=416380
X2670 3143 1 3209 388 2 3217 ND3 $T=540640 507480 1 0 $X=540640 $Y=502060
X2671 3227 1 3241 2913 2 3221 ND3 $T=546220 386520 1 180 $X=543740 $Y=386140
X2672 3263 1 3012 3173 2 3248 ND3 $T=545600 376440 0 0 $X=545600 $Y=376060
X2673 3246 1 3109 3211 2 3239 ND3 $T=548700 386520 0 180 $X=546220 $Y=381100
X2674 3242 1 3250 3251 2 3256 ND3 $T=547460 497400 1 0 $X=547460 $Y=491980
X2675 3231 1 3291 3282 2 3315 ND3 $T=555520 507480 1 0 $X=555520 $Y=502060
X2676 3283 1 3330 3333 2 3089 ND3 $T=559860 487320 0 0 $X=559860 $Y=486940
X2677 3345 1 3341 3033 2 3332 ND3 $T=563580 386520 0 180 $X=561100 $Y=381100
X2678 3404 1 3388 3304 2 3393 ND3 $T=570400 396600 0 0 $X=570400 $Y=396220
X2679 4839 1 4854 746 2 4290 ND3 $T=850640 487320 1 0 $X=850640 $Y=481900
X2680 4853 1 4868 751 2 4523 ND3 $T=853120 487320 1 0 $X=853120 $Y=481900
X2681 4942 1 4936 770 2 4616 ND3 $T=866140 507480 0 180 $X=863660 $Y=502060
X2682 4902 1 5002 798 2 4590 ND3 $T=878540 396600 1 0 $X=878540 $Y=391180
X2683 5025 1 5021 801 2 4705 ND3 $T=884120 517560 0 180 $X=881640 $Y=512140
X2684 5032 1 5029 805 2 4516 ND3 $T=885980 406680 0 180 $X=883500 $Y=401260
X2685 5121 1 5115 813 2 4683 ND3 $T=903340 517560 0 180 $X=900860 $Y=512140
X2686 5188 1 5185 829 2 4546 ND3 $T=915740 517560 0 180 $X=913260 $Y=512140
X2687 20 22 1220 2 1 ND2S $T=225060 537720 0 180 $X=223200 $Y=532300
X2688 1331 1321 1319 2 1 ND2S $T=242420 517560 1 180 $X=240560 $Y=517180
X2689 91 1585 1546 2 1 ND2S $T=293880 366360 1 180 $X=292020 $Y=365980
X2690 1516 1602 1541 2 1 ND2S $T=295740 376440 1 180 $X=293880 $Y=376060
X2691 1509 1598 1558 2 1 ND2S $T=295740 386520 1 180 $X=293880 $Y=386140
X2692 1613 1607 1584 2 1 ND2S $T=300080 396600 0 180 $X=298220 $Y=391180
X2693 1612 1611 1602 2 1 ND2S $T=300700 376440 1 180 $X=298840 $Y=376060
X2694 1579 1640 1560 2 1 ND2S $T=300700 426840 1 180 $X=298840 $Y=426460
X2695 1626 1621 1598 2 1 ND2S $T=301320 386520 0 180 $X=299460 $Y=381100
X2696 1636 1650 1585 2 1 ND2S $T=302560 376440 0 180 $X=300700 $Y=371020
X2697 1631 1641 1627 2 1 ND2S $T=302560 457080 0 180 $X=300700 $Y=451660
X2698 1633 1645 1637 2 1 ND2S $T=302560 406680 0 0 $X=302560 $Y=406300
X2699 1642 1678 1648 2 1 ND2S $T=305040 487320 0 180 $X=303180 $Y=481900
X2700 1675 1670 1641 2 1 ND2S $T=306900 447000 1 180 $X=305040 $Y=446620
X2701 1644 1697 1668 2 1 ND2S $T=308140 386520 1 180 $X=306280 $Y=386140
X2702 1680 1691 1645 2 1 ND2S $T=308140 406680 1 180 $X=306280 $Y=406300
X2703 1686 1657 1599 2 1 ND2S $T=308140 426840 0 180 $X=306280 $Y=421420
X2704 1634 1679 97 2 1 ND2S $T=306900 376440 0 0 $X=306900 $Y=376060
X2705 1646 1711 1706 2 1 ND2S $T=307520 436920 0 0 $X=307520 $Y=436540
X2706 1713 1666 1652 2 1 ND2S $T=310000 416760 1 0 $X=310000 $Y=411340
X2707 1705 1729 1657 2 1 ND2S $T=311860 426840 1 180 $X=310000 $Y=426460
X2708 1699 1730 1649 2 1 ND2S $T=311860 447000 1 180 $X=310000 $Y=446620
X2709 1692 1649 1707 2 1 ND2S $T=310000 467160 1 0 $X=310000 $Y=461740
X2710 1720 1672 1727 2 1 ND2S $T=311240 457080 0 0 $X=311240 $Y=456700
X2711 1704 1738 1666 2 1 ND2S $T=313720 396600 1 180 $X=311860 $Y=396220
X2712 1723 1608 1727 2 1 ND2S $T=311860 426840 1 0 $X=311860 $Y=421420
X2713 1734 1767 1678 2 1 ND2S $T=313720 487320 0 180 $X=311860 $Y=481900
X2714 1660 1752 1607 2 1 ND2S $T=314340 396600 0 180 $X=312480 $Y=391180
X2715 1740 1726 1727 2 1 ND2S $T=314340 467160 1 180 $X=312480 $Y=466780
X2716 1732 1582 1745 2 1 ND2S $T=313100 406680 0 0 $X=313100 $Y=406300
X2717 1733 1698 1745 2 1 ND2S $T=313100 416760 1 0 $X=313100 $Y=411340
X2718 1605 1751 1747 2 1 ND2S $T=313100 497400 1 0 $X=313100 $Y=491980
X2719 1748 1609 1727 2 1 ND2S $T=315580 436920 1 180 $X=313720 $Y=436540
X2720 1756 1743 1727 2 1 ND2S $T=316200 467160 1 180 $X=314340 $Y=466780
X2721 1731 1783 1751 2 1 ND2S $T=316820 497400 0 180 $X=314960 $Y=491980
X2722 1770 1555 111 2 1 ND2S $T=316820 366360 0 0 $X=316820 $Y=365980
X2723 1780 1581 1745 2 1 ND2S $T=316820 386520 1 0 $X=316820 $Y=381100
X2724 1761 1781 1640 2 1 ND2S $T=318680 426840 1 180 $X=316820 $Y=426460
X2725 1731 1715 1784 2 1 ND2S $T=317440 497400 1 0 $X=317440 $Y=491980
X2726 1788 1565 1745 2 1 ND2S $T=318680 396600 1 0 $X=318680 $Y=391180
X2727 1775 1542 1745 2 1 ND2S $T=318680 406680 1 0 $X=318680 $Y=401260
X2728 1784 1808 1778 2 1 ND2S $T=324260 497400 1 0 $X=324260 $Y=491980
X2729 1825 1778 1832 2 1 ND2S $T=327360 497400 1 0 $X=327360 $Y=491980
X2730 1841 1802 1835 2 1 ND2S $T=329840 497400 0 0 $X=329840 $Y=497020
X2731 1881 1875 1835 2 1 ND2S $T=339760 497400 0 0 $X=339760 $Y=497020
X2732 1885 1891 1898 2 1 ND2S $T=341620 517560 1 0 $X=341620 $Y=512140
X2733 1906 1913 1891 2 1 ND2S $T=345960 507480 1 180 $X=344100 $Y=507100
X2734 1922 1918 1815 2 1 ND2S $T=347820 386520 1 180 $X=345960 $Y=386140
X2735 1933 1942 1911 2 1 ND2S $T=350920 376440 1 180 $X=349060 $Y=376060
X2736 1803 1959 1960 2 1 ND2S $T=354020 386520 1 180 $X=352160 $Y=386140
X2737 1906 1975 1998 2 1 ND2S $T=355880 507480 0 0 $X=355880 $Y=507100
X2738 1970 1994 2003 2 1 ND2S $T=359600 517560 1 0 $X=359600 $Y=512140
X2739 155 2011 2033 2 1 ND2S $T=362700 376440 1 0 $X=362700 $Y=371020
X2740 1998 2049 2029 2 1 ND2S $T=366420 507480 0 180 $X=364560 $Y=502060
X2741 2056 2029 2047 2 1 ND2S $T=364560 517560 1 0 $X=364560 $Y=512140
X2742 2100 2083 1835 2 1 ND2S $T=373240 507480 0 180 $X=371380 $Y=502060
X2743 2165 2221 2171 2 1 ND2S $T=386880 507480 0 180 $X=385020 $Y=502060
X2744 2199 2197 2080 2 1 ND2S $T=389360 507480 1 180 $X=387500 $Y=507100
X2745 2213 2220 2221 2 1 ND2S $T=391220 507480 0 0 $X=391220 $Y=507100
X2746 2229 2233 2257 2 1 ND2S $T=393080 517560 1 0 $X=393080 $Y=512140
X2747 2271 2269 2233 2 1 ND2S $T=400520 507480 1 0 $X=400520 $Y=502060
X2748 2283 2278 2080 2 1 ND2S $T=401760 517560 1 0 $X=401760 $Y=512140
X2749 2284 2294 2080 2 1 ND2S $T=405480 507480 1 0 $X=405480 $Y=502060
X2750 2334 2343 203 2 1 ND2S $T=412920 527640 1 180 $X=411060 $Y=527260
X2751 2384 2376 2386 2 1 ND2S $T=419740 497400 0 0 $X=419740 $Y=497020
X2752 2385 2387 2080 2 1 ND2S $T=420980 507480 0 0 $X=420980 $Y=507100
X2753 2403 2391 2386 2 1 ND2S $T=423460 497400 0 0 $X=423460 $Y=497020
X2754 2314 2417 2319 2 1 ND2S $T=425320 507480 0 180 $X=423460 $Y=502060
X2755 2359 2412 2395 2 1 ND2S $T=425940 507480 1 0 $X=425940 $Y=502060
X2756 2440 2426 2414 2 1 ND2S $T=429040 416760 1 180 $X=427180 $Y=416380
X2757 2429 2423 2412 2 1 ND2S $T=429040 497400 0 180 $X=427180 $Y=491980
X2758 2418 2428 2417 2 1 ND2S $T=429660 497400 1 180 $X=427800 $Y=497020
X2759 2418 2456 2429 2 1 ND2S $T=430280 507480 0 0 $X=430280 $Y=507100
X2760 2459 2454 2431 2 1 ND2S $T=434000 517560 0 180 $X=432140 $Y=512140
X2761 2458 2470 2435 2 1 ND2S $T=434000 527640 0 180 $X=432140 $Y=522220
X2762 1921 2463 239 2 1 ND2S $T=434000 396600 0 0 $X=434000 $Y=396220
X2763 2474 2469 236 2 1 ND2S $T=435860 527640 1 180 $X=434000 $Y=527260
X2764 2452 2444 2464 2 1 ND2S $T=435240 426840 1 0 $X=435240 $Y=421420
X2765 2473 2480 2454 2 1 ND2S $T=436480 517560 1 0 $X=436480 $Y=512140
X2766 2511 2504 2470 2 1 ND2S $T=442060 527640 0 180 $X=440200 $Y=522220
X2767 2500 2521 2499 2 1 ND2S $T=444540 457080 0 180 $X=442680 $Y=451660
X2768 2490 2528 2469 2 1 ND2S $T=445160 527640 1 180 $X=443300 $Y=527260
X2769 2569 2568 2560 2 1 ND2S $T=451360 436920 1 180 $X=449500 $Y=436540
X2770 2603 2624 2640 2 1 ND2S $T=461900 457080 1 0 $X=461900 $Y=451660
X2771 2609 2633 2541 2 1 ND2S $T=463760 416760 1 0 $X=463760 $Y=411340
X2772 2592 2640 2625 2 1 ND2S $T=463760 457080 1 0 $X=463760 $Y=451660
X2773 2616 2657 2624 2 1 ND2S $T=466240 436920 0 180 $X=464380 $Y=431500
X2774 2586 2714 2611 2 1 ND2S $T=474920 477240 1 180 $X=473060 $Y=476860
X2775 2702 2703 2642 2 1 ND2S $T=474300 396600 0 0 $X=474300 $Y=396220
X2776 2709 2747 2722 2 1 ND2S $T=478640 447000 0 180 $X=476780 $Y=441580
X2777 2706 2722 2676 2 1 ND2S $T=476780 447000 0 0 $X=476780 $Y=446620
X2778 2674 2764 2747 2 1 ND2S $T=482360 447000 0 180 $X=480500 $Y=441580
X2779 2772 2770 2697 2 1 ND2S $T=484840 376440 1 0 $X=484840 $Y=371020
X2780 2789 2823 2788 2 1 ND2S $T=494140 436920 1 0 $X=494140 $Y=431500
X2781 2809 2853 2849 2 1 ND2S $T=496000 447000 1 0 $X=496000 $Y=441580
X2782 2802 2844 2621 2 1 ND2S $T=496620 406680 0 0 $X=496620 $Y=406300
X2783 2849 2852 2730 2 1 ND2S $T=498480 436920 1 180 $X=496620 $Y=436540
X2784 2875 2871 2621 2 1 ND2S $T=500960 416760 1 180 $X=499100 $Y=416380
X2785 2855 2904 2882 2 1 ND2S $T=505300 436920 0 180 $X=503440 $Y=431500
X2786 2911 2933 2941 2 1 ND2S $T=509020 517560 0 0 $X=509020 $Y=517180
X2787 2928 2926 337 2 1 ND2S $T=509020 527640 0 0 $X=509020 $Y=527260
X2788 2978 2960 340 2 1 ND2S $T=513980 396600 0 180 $X=512120 $Y=391180
X2789 2885 2962 2982 2 1 ND2S $T=512120 497400 0 0 $X=512120 $Y=497020
X2790 2934 2970 327 2 1 ND2S $T=513980 537720 0 180 $X=512120 $Y=532300
X2791 2978 2943 2986 2 1 ND2S $T=512740 396600 0 0 $X=512740 $Y=396220
X2792 2951 2994 2971 2 1 ND2S $T=515220 477240 0 0 $X=515220 $Y=476860
X2793 2826 2995 346 2 1 ND2S $T=515220 497400 0 0 $X=515220 $Y=497020
X2794 2997 2996 2986 2 1 ND2S $T=515840 396600 1 0 $X=515840 $Y=391180
X2795 2997 2923 3008 2 1 ND2S $T=515840 396600 0 0 $X=515840 $Y=396220
X2796 338 2991 351 2 1 ND2S $T=515840 527640 1 0 $X=515840 $Y=522220
X2797 2851 3011 3020 2 1 ND2S $T=517080 497400 0 0 $X=517080 $Y=497020
X2798 348 2963 3025 2 1 ND2S $T=517700 507480 0 0 $X=517700 $Y=507100
X2799 2838 3018 3041 2 1 ND2S $T=519560 487320 0 0 $X=519560 $Y=486940
X2800 321 3019 356 2 1 ND2S $T=519560 507480 1 0 $X=519560 $Y=502060
X2801 2916 3029 3054 2 1 ND2S $T=519560 527640 1 0 $X=519560 $Y=522220
X2802 3033 3043 2948 2 1 ND2S $T=520800 416760 1 0 $X=520800 $Y=411340
X2803 350 3050 3066 2 1 ND2S $T=522660 376440 0 0 $X=522660 $Y=376060
X2804 339 3060 3002 2 1 ND2S $T=524520 416760 0 180 $X=522660 $Y=411340
X2805 2729 3053 3025 2 1 ND2S $T=524520 497400 1 180 $X=522660 $Y=497020
X2806 361 2977 3066 2 1 ND2S $T=523280 366360 0 0 $X=523280 $Y=365980
X2807 3046 3077 365 2 1 ND2S $T=523900 527640 0 0 $X=523900 $Y=527260
X2808 3044 3089 2971 2 1 ND2S $T=524520 467160 1 0 $X=524520 $Y=461740
X2809 2980 3073 2971 2 1 ND2S $T=524520 477240 1 0 $X=524520 $Y=471820
X2810 3084 3118 2919 2 1 ND2S $T=526380 507480 0 180 $X=524520 $Y=502060
X2811 2939 3080 2971 2 1 ND2S $T=525140 457080 0 0 $X=525140 $Y=456700
X2812 2812 3093 2904 2 1 ND2S $T=527000 497400 0 180 $X=525140 $Y=491980
X2813 2909 3085 3095 2 1 ND2S $T=525760 517560 1 0 $X=525760 $Y=512140
X2814 3082 3068 2986 2 1 ND2S $T=528240 406680 0 0 $X=528240 $Y=406300
X2815 3108 3086 3123 2 1 ND2S $T=528860 376440 1 0 $X=528860 $Y=371020
X2816 376 3120 3066 2 1 ND2S $T=531960 386520 0 180 $X=530100 $Y=381100
X2817 3082 3145 340 2 1 ND2S $T=530100 406680 1 0 $X=530100 $Y=401260
X2818 3124 3132 3008 2 1 ND2S $T=530100 406680 0 0 $X=530100 $Y=406300
X2819 3134 3136 321 2 1 ND2S $T=531960 487320 1 180 $X=530100 $Y=486940
X2820 375 3101 3066 2 1 ND2S $T=530720 376440 1 0 $X=530720 $Y=371020
X2821 359 3149 3002 2 1 ND2S $T=532580 416760 0 180 $X=530720 $Y=411340
X2822 3081 3143 321 2 1 ND2S $T=533200 507480 1 180 $X=531340 $Y=507100
X2823 3108 377 3151 2 1 ND2S $T=533200 376440 1 0 $X=533200 $Y=371020
X2824 3158 3155 3008 2 1 ND2S $T=535680 406680 0 180 $X=533820 $Y=401260
X2825 3134 3183 2736 2 1 ND2S $T=536920 487320 0 180 $X=535060 $Y=481900
X2826 3175 3147 2736 2 1 ND2S $T=537540 487320 1 180 $X=535680 $Y=486940
X2827 3150 3138 3154 2 1 ND2S $T=535680 497400 0 0 $X=535680 $Y=497020
X2828 3124 3165 3182 2 1 ND2S $T=536920 406680 0 0 $X=536920 $Y=406300
X2829 3193 3146 2986 2 1 ND2S $T=540640 396600 1 180 $X=538780 $Y=396220
X2830 3175 3196 3154 2 1 ND2S $T=540640 487320 0 180 $X=538780 $Y=481900
X2831 3187 3167 3157 2 1 ND2S $T=539400 366360 0 0 $X=539400 $Y=365980
X2832 3186 3188 3213 2 1 ND2S $T=540640 376440 0 0 $X=540640 $Y=376060
X2833 3078 3189 3182 2 1 ND2S $T=540640 406680 1 0 $X=540640 $Y=401260
X2834 384 3172 3213 2 1 ND2S $T=541260 366360 0 0 $X=541260 $Y=365980
X2835 3187 3178 3213 2 1 ND2S $T=541260 376440 1 0 $X=541260 $Y=371020
X2836 3222 3030 3180 2 1 ND2S $T=543740 416760 1 0 $X=543740 $Y=411340
X2837 3225 389 3157 2 1 ND2S $T=544360 366360 0 0 $X=544360 $Y=365980
X2838 3249 3200 3157 2 1 ND2S $T=544360 376440 1 0 $X=544360 $Y=371020
X2839 3252 3221 3157 2 1 ND2S $T=544360 386520 1 0 $X=544360 $Y=381100
X2840 3237 3227 3182 2 1 ND2S $T=546220 396600 0 180 $X=544360 $Y=391180
X2841 3107 3231 2982 2 1 ND2S $T=544360 507480 1 0 $X=544360 $Y=502060
X2842 3243 3215 3233 2 1 ND2S $T=547460 416760 0 180 $X=545600 $Y=411340
X2843 3222 3181 393 2 1 ND2S $T=546220 406680 0 0 $X=546220 $Y=406300
X2844 3247 3242 3176 2 1 ND2S $T=548080 497400 1 180 $X=546220 $Y=497020
X2845 394 3246 383 2 1 ND2S $T=548700 386520 1 180 $X=546840 $Y=386140
X2846 392 390 3213 2 1 ND2S $T=547460 366360 0 0 $X=547460 $Y=365980
X2847 3238 385 2948 2 1 ND2S $T=548080 396600 0 0 $X=548080 $Y=396220
X2848 397 3263 383 2 1 ND2S $T=549320 376440 0 0 $X=549320 $Y=376060
X2849 3073 3260 3267 2 1 ND2S $T=549320 497400 0 0 $X=549320 $Y=497020
X2850 3205 3250 391 2 1 ND2S $T=549940 497400 1 0 $X=549940 $Y=491980
X2851 371 3277 383 2 1 ND2S $T=553040 386520 0 180 $X=551180 $Y=381100
X2852 3266 3256 3154 2 1 ND2S $T=551180 487320 1 0 $X=551180 $Y=481900
X2853 3175 3283 3281 2 1 ND2S $T=554280 497400 0 180 $X=552420 $Y=491980
X2854 394 3264 393 2 1 ND2S $T=553040 386520 1 0 $X=553040 $Y=381100
X2855 3205 3291 374 2 1 ND2S $T=553660 507480 1 0 $X=553660 $Y=502060
X2856 3247 3293 3268 2 1 ND2S $T=554280 497400 0 0 $X=554280 $Y=497020
X2857 3229 3307 3279 2 1 ND2S $T=556760 426840 1 180 $X=554900 $Y=426460
X2858 3286 3279 3312 2 1 ND2S $T=554900 436920 1 0 $X=554900 $Y=431500
X2859 3261 3312 3254 2 1 ND2S $T=556760 436920 1 180 $X=554900 $Y=436540
X2860 3205 3300 401 2 1 ND2S $T=556760 497400 0 180 $X=554900 $Y=491980
X2861 3247 3315 3271 2 1 ND2S $T=558000 507480 1 0 $X=558000 $Y=502060
X2862 3336 3332 3346 2 1 ND2S $T=561720 386520 0 0 $X=561720 $Y=386140
X2863 3344 3303 3354 2 1 ND2S $T=562960 366360 0 0 $X=562960 $Y=365980
X2864 3297 3133 411 2 1 ND2S $T=564200 386520 0 0 $X=564200 $Y=386140
X2865 3362 3272 3370 2 1 ND2S $T=566060 406680 1 0 $X=566060 $Y=401260
X2866 417 3345 3360 2 1 ND2S $T=569780 386520 1 0 $X=569780 $Y=381100
X2867 3424 3405 427 2 1 ND2S $T=574120 376440 1 0 $X=574120 $Y=371020
X2868 3395 3414 3422 2 1 ND2S $T=575980 436920 0 0 $X=575980 $Y=436540
X2869 3398 3422 3364 2 1 ND2S $T=577840 447000 0 180 $X=575980 $Y=441580
X2870 3476 3455 3442 2 1 ND2S $T=583420 376440 0 0 $X=583420 $Y=376060
X2871 3471 3466 3476 2 1 ND2S $T=585280 386520 1 0 $X=585280 $Y=381100
X2872 446 3442 448 2 1 ND2S $T=587140 376440 1 0 $X=587140 $Y=371020
X2873 3509 3496 3520 2 1 ND2S $T=590240 386520 0 0 $X=590240 $Y=386140
X2874 3510 3500 3521 2 1 ND2S $T=590240 406680 0 0 $X=590240 $Y=406300
X2875 3510 3512 3525 2 1 ND2S $T=590860 416760 1 0 $X=590860 $Y=411340
X2876 3510 3501 3522 2 1 ND2S $T=590860 416760 0 0 $X=590860 $Y=416380
X2877 3523 3520 451 2 1 ND2S $T=593340 386520 0 180 $X=591480 $Y=381100
X2878 3532 3452 3537 2 1 ND2S $T=593960 426840 1 0 $X=593960 $Y=421420
X2879 3528 3497 3548 2 1 ND2S $T=595820 396600 1 0 $X=595820 $Y=391180
X2880 3470 3538 3473 2 1 ND2S $T=595820 447000 0 0 $X=595820 $Y=446620
X2881 3518 3550 3558 2 1 ND2S $T=597680 517560 1 0 $X=597680 $Y=512140
X2882 3522 3498 3568 2 1 ND2S $T=598300 426840 1 0 $X=598300 $Y=421420
X2883 3532 3579 3569 2 1 ND2S $T=598920 426840 0 0 $X=598920 $Y=426460
X2884 3565 3548 3560 2 1 ND2S $T=602020 396600 0 180 $X=600160 $Y=391180
X2885 3573 3477 3580 2 1 ND2S $T=600780 416760 1 0 $X=600780 $Y=411340
X2886 3583 3580 3593 2 1 ND2S $T=602640 396600 0 0 $X=602640 $Y=396220
X2887 3569 3516 3606 2 1 ND2S $T=605120 436920 1 0 $X=605120 $Y=431500
X2888 3567 3469 3613 2 1 ND2S $T=605740 416760 0 0 $X=605740 $Y=416380
X2889 3642 3613 3635 2 1 ND2S $T=611320 416760 0 0 $X=611320 $Y=416380
X2890 3669 3600 3651 2 1 ND2S $T=612560 436920 0 0 $X=612560 $Y=436540
X2891 3678 3568 3664 2 1 ND2S $T=613800 426840 1 0 $X=613800 $Y=421420
X2892 3673 3672 3684 2 1 ND2S $T=615040 447000 1 0 $X=615040 $Y=441580
X2893 3665 3603 3686 2 1 ND2S $T=615660 426840 0 0 $X=615660 $Y=426460
X2894 3829 3854 3839 2 1 ND2S $T=647280 507480 0 180 $X=645420 $Y=502060
X2895 3815 3888 3741 2 1 ND2S $T=649760 477240 0 0 $X=649760 $Y=476860
X2896 4101 4100 4037 2 1 ND2S $T=690060 497400 1 180 $X=688200 $Y=497020
X2897 4088 4081 4018 2 1 ND2S $T=690060 507480 1 180 $X=688200 $Y=507100
X2898 4116 4115 4038 2 1 ND2S $T=693780 447000 1 180 $X=691920 $Y=446620
X2899 4139 4121 4048 2 1 ND2S $T=696880 426840 1 180 $X=695020 $Y=426460
X2900 4135 4134 4057 2 1 ND2S $T=697500 436920 1 180 $X=695640 $Y=436540
X2901 4165 4149 563 2 1 ND2S $T=702460 537720 0 180 $X=700600 $Y=532300
X2902 4151 4194 4016 2 1 ND2S $T=708040 497400 1 180 $X=706180 $Y=497020
X2903 4253 4284 4291 2 1 ND2S $T=727260 436920 1 0 $X=727260 $Y=431500
X2904 4317 4298 4289 2 1 ND2S $T=732840 436920 0 180 $X=730980 $Y=431500
X2905 5504 5483 5503 2 1 ND2S $T=987040 467160 1 0 $X=987040 $Y=461740
X2906 5585 5578 5580 2 1 ND2S $T=1003780 376440 0 180 $X=1001920 $Y=371020
X2907 5581 5535 5589 2 1 ND2S $T=1002540 467160 0 0 $X=1002540 $Y=466780
X2908 5700 5518 5708 2 1 ND2S $T=1027960 376440 1 0 $X=1027960 $Y=371020
X2909 1036 5450 5715 2 1 ND2S $T=1029200 366360 0 0 $X=1029200 $Y=365980
X2910 5720 5583 5730 2 1 ND2S $T=1032300 467160 0 0 $X=1032300 $Y=466780
X2911 5827 5506 5823 2 1 ND2S $T=1052140 467160 0 0 $X=1052140 $Y=466780
X2912 1242 20 1 5 1228 1223 2 MOAI1S $T=226920 517560 1 180 $X=223200 $Y=517180
X2913 2680 285 1 2475 2652 2692 2 MOAI1S $T=469340 416760 1 0 $X=469340 $Y=411340
X2914 1982 2680 1 2475 2730 2755 2 MOAI1S $T=476160 406680 1 0 $X=476160 $Y=401260
X2915 2680 2463 1 2475 2734 2732 2 MOAI1S $T=476780 396600 1 0 $X=476780 $Y=391180
X2916 1936 2680 1 2475 2753 2744 2 MOAI1S $T=479260 416760 1 0 $X=479260 $Y=411340
X2917 2793 2799 1 2793 2799 2817 2 MOAI1S $T=489180 426840 0 0 $X=489180 $Y=426460
X2918 2809 2705 1 2809 2705 2827 2 MOAI1S $T=491660 416760 1 0 $X=491660 $Y=411340
X2919 2838 2667 1 2723 2695 2846 2 MOAI1S $T=500340 487320 1 180 $X=496620 $Y=486940
X2920 2843 2869 1 2861 240 2854 2 MOAI1S $T=501580 406680 0 180 $X=497860 $Y=401260
X2921 2851 2839 1 2723 2737 2859 2 MOAI1S $T=501580 497400 0 180 $X=497860 $Y=491980
X2922 2821 2869 1 2861 2533 2856 2 MOAI1S $T=502200 406680 1 180 $X=498480 $Y=406300
X2923 2834 2730 1 2834 2730 2882 2 MOAI1S $T=499100 436920 1 0 $X=499100 $Y=431500
X2924 2826 2857 1 2867 2746 2877 2 MOAI1S $T=499100 497400 0 0 $X=499100 $Y=497020
X2925 2885 2839 1 2890 2723 2912 2 MOAI1S $T=502820 497400 1 0 $X=502820 $Y=491980
X2926 2792 2869 1 2906 2421 2908 2 MOAI1S $T=504060 426840 0 0 $X=504060 $Y=426460
X2927 2916 2857 1 2867 2899 2898 2 MOAI1S $T=507780 507480 0 180 $X=504060 $Y=502060
X2928 338 2857 1 2867 2891 2896 2 MOAI1S $T=507780 517560 1 180 $X=504060 $Y=517180
X2929 2874 2914 1 2905 329 2900 2 MOAI1S $T=508400 386520 0 180 $X=504680 $Y=381100
X2930 2833 2884 1 2906 2687 2939 2 MOAI1S $T=507780 426840 0 0 $X=507780 $Y=426460
X2931 2883 2914 1 2905 323 2945 2 MOAI1S $T=509020 376440 0 0 $X=509020 $Y=376060
X2932 334 2914 1 2905 2420 2922 2 MOAI1S $T=512740 386520 1 180 $X=509020 $Y=386140
X2933 345 2884 1 2906 2530 2949 2 MOAI1S $T=515220 426840 1 180 $X=511500 $Y=426460
X2934 342 2914 1 2905 223 2998 2 MOAI1S $T=512740 386520 1 0 $X=512740 $Y=381100
X2935 332 2884 1 2989 2556 2967 2 MOAI1S $T=518320 436920 0 180 $X=514600 $Y=431500
X2936 2667 2966 1 2866 3009 3010 2 MOAI1S $T=514600 436920 0 0 $X=514600 $Y=436540
X2937 348 2857 1 347 2867 2975 2 MOAI1S $T=519560 517560 0 180 $X=515840 $Y=512140
X2938 331 2914 1 2905 358 3035 2 MOAI1S $T=518940 396600 1 0 $X=518940 $Y=391180
X2939 3006 108 1 2866 3038 3031 2 MOAI1S $T=518940 447000 1 0 $X=518940 $Y=441580
X2940 2667 2664 1 2866 3047 3051 2 MOAI1S $T=519560 436920 0 0 $X=519560 $Y=436540
X2941 2974 2914 1 2906 362 3061 2 MOAI1S $T=520800 426840 0 0 $X=520800 $Y=426460
X2942 2909 2857 1 2867 363 3039 2 MOAI1S $T=521420 517560 0 0 $X=521420 $Y=517180
X2943 3046 2857 1 2867 364 3065 2 MOAI1S $T=522040 517560 1 0 $X=522040 $Y=512140
X2944 3081 372 1 3093 3053 3084 2 MOAI1S $T=529480 507480 1 180 $X=525760 $Y=507100
X2945 3094 2884 1 2906 3115 3128 2 MOAI1S $T=527000 436920 1 0 $X=527000 $Y=431500
X2946 3064 3204 1 3119 3244 3218 2 MOAI1S $T=544360 487320 1 0 $X=544360 $Y=481900
X2947 3967 3955 1 3967 3971 3958 2 MOAI1S $T=667120 497400 1 180 $X=663400 $Y=497020
X2948 523 3656 1 523 3971 3965 2 MOAI1S $T=675800 497400 0 180 $X=672080 $Y=491980
X2949 4019 3736 1 4019 535 4011 2 MOAI1S $T=677660 527640 1 180 $X=673940 $Y=527260
X2950 4019 3820 1 4019 3971 4023 2 MOAI1S $T=683240 497400 0 180 $X=679520 $Y=491980
X2951 4053 3703 1 4053 545 4006 2 MOAI1S $T=686960 517560 0 180 $X=683240 $Y=512140
X2952 4077 4034 1 4077 4073 4084 2 MOAI1S $T=685720 497400 1 0 $X=685720 $Y=491980
X2953 4089 4017 1 4089 4087 4005 2 MOAI1S $T=691920 447000 0 180 $X=688200 $Y=441580
X2954 4099 4050 1 4099 549 4031 2 MOAI1S $T=693160 487320 0 180 $X=689440 $Y=481900
X2955 4105 4068 1 4105 4103 4028 2 MOAI1S $T=693780 426840 0 180 $X=690060 $Y=421420
X2956 4105 4029 1 4105 4087 4083 2 MOAI1S $T=695640 447000 0 180 $X=691920 $Y=441580
X2957 4077 4063 1 4077 554 4086 2 MOAI1S $T=695640 497400 1 180 $X=691920 $Y=497020
X2958 4118 4130 1 4118 554 4082 2 MOAI1S $T=697500 406680 0 180 $X=693780 $Y=401260
X2959 4118 4117 1 4118 4087 4055 2 MOAI1S $T=697500 416760 1 180 $X=693780 $Y=416380
X2960 4089 3960 1 4089 4103 4035 2 MOAI1S $T=697500 436920 0 180 $X=693780 $Y=431500
X2961 4119 3851 1 4119 549 4049 2 MOAI1S $T=697500 477240 0 180 $X=693780 $Y=471820
X2962 4119 4126 1 4119 4073 4157 2 MOAI1S $T=695020 457080 0 0 $X=695020 $Y=456700
X2963 4120 4127 1 4120 545 4145 2 MOAI1S $T=695020 507480 0 0 $X=695020 $Y=507100
X2964 4146 4153 1 4146 4087 4078 2 MOAI1S $T=701220 416760 0 180 $X=697500 $Y=411340
X2965 4146 4125 1 4146 554 4067 2 MOAI1S $T=702460 396600 1 180 $X=698740 $Y=396220
X2966 4019 4085 1 4019 554 4162 2 MOAI1S $T=698740 497400 1 0 $X=698740 $Y=491980
X2967 4118 4168 1 4118 4103 4186 2 MOAI1S $T=701840 406680 1 0 $X=701840 $Y=401260
X2968 4146 4047 1 4146 4103 4164 2 MOAI1S $T=705560 416760 0 180 $X=701840 $Y=411340
X2969 4172 4102 1 4172 4087 4094 2 MOAI1S $T=706180 396600 0 180 $X=702460 $Y=391180
X2970 4173 570 1 4173 549 565 2 MOAI1S $T=706180 537720 0 180 $X=702460 $Y=532300
X2971 4120 3735 1 4120 4179 4185 2 MOAI1S $T=703700 507480 0 0 $X=703700 $Y=507100
X2972 4172 4075 1 4172 4103 4108 2 MOAI1S $T=708040 386520 1 180 $X=704320 $Y=386140
X2973 4077 4178 1 4077 4179 4198 2 MOAI1S $T=704940 507480 1 0 $X=704940 $Y=502060
X2974 4099 4181 1 4188 4073 4193 2 MOAI1S $T=705560 467160 0 0 $X=705560 $Y=466780
X2975 4192 4196 1 4192 4087 4183 2 MOAI1S $T=710520 396600 0 180 $X=706800 $Y=391180
X2976 4053 3838 1 4053 566 4180 2 MOAI1S $T=710520 517560 0 180 $X=706800 $Y=512140
X2977 4192 4163 1 4192 4103 4158 2 MOAI1S $T=711760 376440 1 180 $X=708040 $Y=376060
X2978 4099 3797 1 4099 4179 4207 2 MOAI1S $T=709280 467160 0 0 $X=709280 $Y=466780
X2979 4119 4213 1 4205 4179 4201 2 MOAI1S $T=714240 477240 0 180 $X=710520 $Y=471820
X2980 4197 3869 1 4197 4179 4175 2 MOAI1S $T=714240 497400 0 180 $X=710520 $Y=491980
X2981 582 3842 1 4053 578 576 2 MOAI1S $T=714240 537720 0 180 $X=710520 $Y=532300
X2982 4022 3824 1 4022 4073 4174 2 MOAI1S $T=716720 447000 0 0 $X=716720 $Y=446620
X2983 4220 3979 1 4036 4073 4233 2 MOAI1S $T=716720 457080 0 0 $X=716720 $Y=456700
X2984 4210 4258 1 4210 4263 4259 2 MOAI1S $T=727260 436920 0 180 $X=723540 $Y=431500
X2985 4268 4283 1 4268 4263 4250 2 MOAI1S $T=729120 426840 1 180 $X=725400 $Y=426460
X2986 4215 594 1 4215 4263 597 2 MOAI1S $T=731600 386520 1 0 $X=731600 $Y=381100
X2987 4231 4044 1 4231 4263 4330 2 MOAI1S $T=732840 426840 1 0 $X=732840 $Y=421420
X2988 4322 4328 1 4322 4263 4347 2 MOAI1S $T=734700 386520 0 0 $X=734700 $Y=386140
X2989 4356 610 1 4239 4263 4286 2 MOAI1S $T=744000 396600 1 180 $X=740280 $Y=396220
X2990 4728 702 1 4754 4757 4724 2 MOAI1S $T=828940 426840 0 0 $X=828940 $Y=426460
X2991 4752 4765 1 4752 4757 4748 2 MOAI1S $T=835140 447000 0 180 $X=831420 $Y=441580
X2992 4752 4767 1 4752 704 4740 2 MOAI1S $T=835140 467160 0 180 $X=831420 $Y=461740
X2993 4776 717 1 4776 704 4726 2 MOAI1S $T=838860 447000 0 180 $X=835140 $Y=441580
X2994 4805 720 1 4779 4757 4786 2 MOAI1S $T=840100 426840 1 180 $X=836380 $Y=426460
X2995 4776 4811 1 4776 4757 4803 2 MOAI1S $T=843200 447000 0 180 $X=839480 $Y=441580
X2996 4822 733 1 4822 4757 4789 2 MOAI1S $T=846920 447000 0 180 $X=843200 $Y=441580
X2997 4820 4833 1 4820 4757 4847 2 MOAI1S $T=847540 447000 0 0 $X=847540 $Y=446620
X2998 4928 778 1 4928 4970 4973 2 MOAI1S $T=869240 426840 0 0 $X=869240 $Y=426460
X2999 4898 4975 1 4898 777 4925 2 MOAI1S $T=874200 447000 1 180 $X=870480 $Y=446620
X3000 4926 4968 1 4926 777 4977 2 MOAI1S $T=871100 467160 1 0 $X=871100 $Y=461740
X3001 4958 4980 1 4958 4970 5000 2 MOAI1S $T=874200 436920 1 0 $X=874200 $Y=431500
X3002 4830 5095 1 4830 704 5074 2 MOAI1S $T=899000 426840 1 180 $X=895280 $Y=426460
X3003 4805 5114 1 4805 704 5079 2 MOAI1S $T=903340 426840 1 180 $X=899620 $Y=426460
X3004 5092 5109 1 5092 819 5052 2 MOAI1S $T=900860 467160 1 0 $X=900860 $Y=461740
X3005 5027 818 1 5027 5133 5061 2 MOAI1S $T=902720 457080 0 0 $X=902720 $Y=456700
X3006 5127 823 1 5127 5125 5068 2 MOAI1S $T=907060 447000 0 180 $X=903340 $Y=441580
X3007 5138 5150 1 5138 5125 5064 2 MOAI1S $T=908920 457080 0 180 $X=905200 $Y=451660
X3008 5127 5162 1 5127 825 5106 2 MOAI1S $T=911400 447000 0 180 $X=907680 $Y=441580
X3009 4923 5157 1 4923 5167 5160 2 MOAI1S $T=908300 426840 0 0 $X=908300 $Y=426460
X3010 5138 5168 1 5138 830 5206 2 MOAI1S $T=911400 467160 1 0 $X=911400 $Y=461740
X3011 5092 5189 1 5092 5133 5200 2 MOAI1S $T=915120 457080 0 0 $X=915120 $Y=456700
X3012 4886 5191 1 4886 5167 5214 2 MOAI1S $T=915740 426840 0 0 $X=915740 $Y=426460
X3013 5138 5136 1 5138 825 5209 2 MOAI1S $T=915740 447000 0 0 $X=915740 $Y=446620
X3014 4830 840 1 4830 5167 5159 2 MOAI1S $T=920700 416760 0 180 $X=916980 $Y=411340
X3015 5192 5172 1 5192 5219 5216 2 MOAI1S $T=918840 497400 1 0 $X=918840 $Y=491980
X3016 5192 5210 1 5192 5133 5223 2 MOAI1S $T=919460 457080 0 0 $X=919460 $Y=456700
X3017 5222 845 1 5222 844 5215 2 MOAI1S $T=925040 386520 1 180 $X=921320 $Y=386140
X3018 4805 5232 1 4805 5167 5218 2 MOAI1S $T=925040 416760 0 180 $X=921320 $Y=411340
X3019 5126 5238 1 5126 5219 5229 2 MOAI1S $T=926280 497400 0 180 $X=922560 $Y=491980
X3020 5235 5239 1 5235 844 5250 2 MOAI1S $T=925040 386520 1 0 $X=925040 $Y=381100
X3021 5241 5253 1 5241 825 5228 2 MOAI1S $T=929380 447000 0 180 $X=925660 $Y=441580
X3022 5241 851 1 5241 5125 5220 2 MOAI1S $T=930620 457080 1 180 $X=926900 $Y=456700
X3023 5222 852 1 5222 819 5245 2 MOAI1S $T=931240 386520 1 180 $X=927520 $Y=386140
X3024 5265 855 1 5265 5133 5277 2 MOAI1S $T=930620 477240 1 0 $X=930620 $Y=471820
X3025 5265 862 1 5265 825 5288 2 MOAI1S $T=933100 447000 1 0 $X=933100 $Y=441580
X3026 5235 5279 1 5235 819 5294 2 MOAI1S $T=933720 386520 1 0 $X=933720 $Y=381100
X3027 5122 866 1 5122 819 5306 2 MOAI1S $T=934340 406680 0 0 $X=934340 $Y=406300
X3028 5292 5300 1 5292 5167 5276 2 MOAI1S $T=939920 416760 1 180 $X=936200 $Y=416380
X3029 5222 875 1 5222 877 5319 2 MOAI1S $T=938680 396600 1 0 $X=938680 $Y=391180
X3030 5265 5304 1 5265 5125 5317 2 MOAI1S $T=938680 457080 1 0 $X=938680 $Y=451660
X3031 5212 5312 1 5212 5167 5334 2 MOAI1S $T=940540 416760 0 0 $X=940540 $Y=416380
X3032 5235 5313 1 5235 877 5330 2 MOAI1S $T=941160 386520 1 0 $X=941160 $Y=381100
X3033 4951 5322 1 4951 877 884 2 MOAI1S $T=943020 366360 0 0 $X=943020 $Y=365980
X3034 5048 881 1 5048 5219 5336 2 MOAI1S $T=943640 497400 1 0 $X=943640 $Y=491980
X3035 5332 889 1 5332 5320 5293 2 MOAI1S $T=948600 447000 1 180 $X=944880 $Y=446620
X3036 5338 896 1 5338 5320 5337 2 MOAI1S $T=951080 436920 0 180 $X=947360 $Y=431500
X3037 5338 5350 1 5338 5125 5325 2 MOAI1S $T=951080 467160 0 180 $X=947360 $Y=461740
X3038 5104 5356 1 5104 5219 5373 2 MOAI1S $T=951080 487320 0 0 $X=951080 $Y=486940
X3039 5332 5368 1 5332 5125 5342 2 MOAI1S $T=955420 467160 0 180 $X=951700 $Y=461740
X3040 5292 907 1 5292 5320 5347 2 MOAI1S $T=957280 396600 0 180 $X=953560 $Y=391180
X3041 5363 5212 1 5212 5320 5380 2 MOAI1S $T=953560 406680 0 0 $X=953560 $Y=406300
X3042 5366 5369 1 5369 909 5383 2 MOAI1S $T=954180 386520 0 0 $X=954180 $Y=386140
X3043 908 912 1 912 909 5391 2 MOAI1S $T=956660 366360 0 0 $X=956660 $Y=365980
X3044 5369 915 1 5369 5327 5394 2 MOAI1S $T=957280 396600 1 0 $X=957280 $Y=391180
X3045 5259 916 1 5259 5393 5397 2 MOAI1S $T=957280 497400 1 0 $X=957280 $Y=491980
X3046 5321 5396 1 5321 5393 5409 2 MOAI1S $T=959760 487320 0 0 $X=959760 $Y=486940
X3047 5402 5405 1 5402 5413 5417 2 MOAI1S $T=961620 477240 1 0 $X=961620 $Y=471820
X3048 5292 922 1 5292 5327 5419 2 MOAI1S $T=962860 406680 0 0 $X=962860 $Y=406300
X3049 5402 5407 1 5402 5416 5420 2 MOAI1S $T=962860 447000 1 0 $X=962860 $Y=441580
X3050 5403 5421 1 5403 5413 5428 2 MOAI1S $T=965340 477240 0 0 $X=965340 $Y=476860
X3051 5403 5425 1 5403 5416 5433 2 MOAI1S $T=966580 447000 1 0 $X=966580 $Y=441580
X3052 5402 5431 1 5402 5378 5426 2 MOAI1S $T=970920 457080 0 180 $X=967200 $Y=451660
X3053 5442 930 1 5442 5327 5439 2 MOAI1S $T=975880 436920 0 180 $X=972160 $Y=431500
X3054 5444 5447 1 5444 924 5390 2 MOAI1S $T=976500 416760 1 180 $X=972780 $Y=416380
X3055 5444 5443 1 5444 5327 5438 2 MOAI1S $T=977740 426840 0 180 $X=974020 $Y=421420
X3056 932 937 1 932 931 5418 2 MOAI1S $T=977740 527640 0 180 $X=974020 $Y=522220
X3057 5403 933 1 5403 5378 5458 2 MOAI1S $T=974640 467160 1 0 $X=974640 $Y=461740
X3058 5442 5465 1 5442 924 5411 2 MOAI1S $T=980220 416760 0 180 $X=976500 $Y=411340
X3059 5454 5459 1 5454 5413 5423 2 MOAI1S $T=980220 507480 1 180 $X=976500 $Y=507100
X3060 5467 5474 1 5467 5413 5453 2 MOAI1S $T=982080 497400 1 180 $X=978360 $Y=497020
X3061 932 948 1 932 944 5415 2 MOAI1S $T=982080 527640 1 180 $X=978360 $Y=527260
X3062 5468 949 1 5468 946 5422 2 MOAI1S $T=982700 376440 1 180 $X=978980 $Y=376060
X3063 5475 952 1 5475 924 5432 2 MOAI1S $T=983320 396600 0 180 $X=979600 $Y=391180
X3064 5454 5494 1 5454 931 5482 2 MOAI1S $T=986420 507480 1 180 $X=982700 $Y=507100
X3065 958 961 1 958 944 5473 2 MOAI1S $T=986420 527640 1 180 $X=982700 $Y=527260
X3066 5489 963 1 5489 5413 5469 2 MOAI1S $T=987040 487320 1 180 $X=983320 $Y=486940
X3067 5500 5509 1 5500 5413 5487 2 MOAI1S $T=988900 477240 0 180 $X=985180 $Y=471820
X3068 5468 966 1 5468 960 5476 2 MOAI1S $T=989520 376440 0 180 $X=985800 $Y=371020
X3069 5475 5521 1 5475 946 5507 2 MOAI1S $T=991380 386520 1 180 $X=987660 $Y=386140
X3070 5511 5522 1 5511 5416 5485 2 MOAI1S $T=991380 426840 1 180 $X=987660 $Y=426460
X3071 5475 971 1 5475 976 5531 2 MOAI1S $T=988280 396600 1 0 $X=988280 $Y=391180
X3072 5454 5529 1 5454 970 5470 2 MOAI1S $T=992000 517560 0 180 $X=988280 $Y=512140
X3073 5527 5533 1 5527 864 5513 2 MOAI1S $T=993240 467160 0 180 $X=989520 $Y=461740
X3074 5467 5534 1 5467 931 5536 2 MOAI1S $T=991380 507480 0 0 $X=991380 $Y=507100
X3075 958 983 1 958 931 5544 2 MOAI1S $T=997580 527640 1 180 $X=993860 $Y=527260
X3076 5549 5514 1 5549 5416 5562 2 MOAI1S $T=995720 436920 1 0 $X=995720 $Y=431500
X3077 5489 5561 1 5489 970 5539 2 MOAI1S $T=999440 487320 1 180 $X=995720 $Y=486940
X3078 5560 5565 1 5560 864 5572 2 MOAI1S $T=998820 457080 0 0 $X=998820 $Y=456700
X3079 5570 5576 1 5570 970 5546 2 MOAI1S $T=1002540 507480 1 180 $X=998820 $Y=507100
X3080 5500 5569 1 5500 5579 5584 2 MOAI1S $T=999440 477240 1 0 $X=999440 $Y=471820
X3081 5468 998 1 5468 976 5550 2 MOAI1S $T=1006880 386520 1 180 $X=1003160 $Y=386140
X3082 5527 5592 1 5527 5579 5622 2 MOAI1S $T=1003780 477240 1 0 $X=1003780 $Y=471820
X3083 5549 5600 1 5549 5588 5575 2 MOAI1S $T=1008120 436920 0 180 $X=1004400 $Y=431500
X3084 5457 5616 1 5457 5579 5597 2 MOAI1S $T=1008120 447000 1 180 $X=1004400 $Y=446620
X3085 5604 5617 1 5604 5601 5598 2 MOAI1S $T=1008120 497400 0 180 $X=1004400 $Y=491980
X3086 5560 5608 1 5560 5579 5619 2 MOAI1S $T=1005020 457080 0 0 $X=1005020 $Y=456700
X3087 5596 5621 1 5596 5588 5635 2 MOAI1S $T=1006880 386520 0 0 $X=1006880 $Y=386140
X3088 5603 5626 1 5603 5588 5636 2 MOAI1S $T=1007500 426840 1 0 $X=1007500 $Y=421420
X3089 5466 5637 1 5466 5579 5627 2 MOAI1S $T=1011840 447000 1 180 $X=1008120 $Y=446620
X3090 5571 5631 1 5571 5588 5643 2 MOAI1S $T=1009360 406680 0 0 $X=1009360 $Y=406300
X3091 5640 1011 1 5640 5588 5654 2 MOAI1S $T=1011220 386520 0 0 $X=1011220 $Y=386140
X3092 5644 5645 1 5644 5652 5657 2 MOAI1S $T=1012460 497400 1 0 $X=1012460 $Y=491980
X3093 5570 5632 1 5570 1005 5620 2 MOAI1S $T=1017420 507480 1 180 $X=1013700 $Y=507100
X3094 5615 5649 1 5615 5588 5661 2 MOAI1S $T=1014320 426840 0 0 $X=1014320 $Y=426460
X3095 1015 5655 1 1015 1016 5665 2 MOAI1S $T=1014940 527640 0 0 $X=1014940 $Y=527260
X3096 5658 1017 1 5658 5652 5630 2 MOAI1S $T=1019280 477240 1 180 $X=1015560 $Y=476860
X3097 5570 1018 1 5570 1021 5673 2 MOAI1S $T=1017420 507480 0 0 $X=1017420 $Y=507100
X3098 5642 1026 1 5642 1005 5684 2 MOAI1S $T=1022380 517560 1 0 $X=1022380 $Y=512140
X3099 5699 5697 1 5560 5652 5677 2 MOAI1S $T=1027340 467160 1 180 $X=1023620 $Y=466780
X3100 5687 1032 1 5687 5601 5667 2 MOAI1S $T=1027340 497400 0 180 $X=1023620 $Y=491980
X3101 5457 1038 1 5681 5652 5689 2 MOAI1S $T=1029200 447000 1 0 $X=1029200 $Y=441580
X3102 1037 5653 1 1037 1016 5721 2 MOAI1S $T=1029200 537720 1 0 $X=1029200 $Y=532300
X3103 5644 5724 1 5644 1021 5734 2 MOAI1S $T=1031060 507480 0 0 $X=1031060 $Y=507100
X3104 1044 5737 1 1044 1016 5744 2 MOAI1S $T=1034160 537720 1 0 $X=1034160 $Y=532300
X3105 5642 1049 1 5642 5742 5763 2 MOAI1S $T=1036640 517560 1 0 $X=1036640 $Y=512140
X3106 5761 5767 1 5761 5742 5750 2 MOAI1S $T=1042840 426840 1 180 $X=1039120 $Y=426460
X3107 5687 1051 1 5687 5742 5770 2 MOAI1S $T=1039120 497400 0 0 $X=1039120 $Y=497020
X3108 5768 5745 1 5768 5652 5783 2 MOAI1S $T=1042220 447000 1 0 $X=1042220 $Y=441580
X3109 5771 5769 1 5771 5652 5781 2 MOAI1S $T=1043460 467160 0 0 $X=1043460 $Y=466780
X3110 5771 1064 1 5771 5601 5796 2 MOAI1S $T=1051520 467160 1 180 $X=1047800 $Y=466780
X3111 5768 5819 1 5768 5601 5812 2 MOAI1S $T=1054000 447000 0 180 $X=1050280 $Y=441580
X3112 5699 1079 1 5699 5601 5861 2 MOAI1S $T=1059580 477240 1 0 $X=1059580 $Y=471820
X3113 5681 5857 1 5681 5601 5872 2 MOAI1S $T=1060200 447000 0 0 $X=1060200 $Y=446620
X3114 1546 2 1591 91 1 NR2 $T=292020 376440 1 0 $X=292020 $Y=371020
X3115 1541 2 1590 1516 1 NR2 $T=293880 386520 1 0 $X=293880 $Y=381100
X3116 1558 2 1610 1509 1 NR2 $T=293880 396600 1 0 $X=293880 $Y=391180
X3117 1584 2 1635 1613 1 NR2 $T=299460 406680 1 0 $X=299460 $Y=401260
X3118 1627 2 1629 1631 1 NR2 $T=300700 447000 0 0 $X=300700 $Y=446620
X3119 1591 2 1634 1590 1 NR2 $T=303180 386520 0 180 $X=301320 $Y=381100
X3120 1610 2 1644 1635 1 NR2 $T=301320 396600 1 0 $X=301320 $Y=391180
X3121 1637 2 1667 1633 1 NR2 $T=304420 406680 0 180 $X=302560 $Y=401260
X3122 1689 2 1668 1667 1 NR2 $T=308140 396600 1 180 $X=306280 $Y=396220
X3123 1599 2 1638 1686 1 NR2 $T=306280 426840 0 0 $X=306280 $Y=426460
X3124 1679 2 1701 1697 1 NR2 $T=306900 386520 1 0 $X=306900 $Y=381100
X3125 1648 2 1694 1642 1 NR2 $T=308140 487320 0 0 $X=308140 $Y=486940
X3126 1694 2 1683 1715 1 NR2 $T=308140 497400 1 0 $X=308140 $Y=491980
X3127 1712 2 1706 1629 1 NR2 $T=311240 447000 0 180 $X=309380 $Y=441580
X3128 1707 2 1712 1692 1 NR2 $T=311240 457080 1 180 $X=309380 $Y=456700
X3129 1652 2 1689 1713 1 NR2 $T=311860 406680 1 180 $X=310000 $Y=406300
X3130 1747 2 1759 1605 1 NR2 $T=314960 497400 1 180 $X=313100 $Y=497020
X3131 1832 2 1797 1825 1 NR2 $T=329220 497400 1 180 $X=327360 $Y=497020
X3132 1888 2 1882 129 1 NR2 $T=341620 376440 1 180 $X=339760 $Y=376060
X3133 1796 2 1886 1862 1 NR2 $T=340380 386520 0 0 $X=340380 $Y=386140
X3134 1844 2 1888 1892 1 NR2 $T=341620 376440 1 0 $X=341620 $Y=371020
X3135 1721 2 1892 1894 1 NR2 $T=341620 376440 0 0 $X=341620 $Y=376060
X3136 1844 2 1915 1721 1 NR2 $T=344100 376440 1 0 $X=344100 $Y=371020
X3137 1967 2 1958 1972 1 NR2 $T=352780 457080 0 0 $X=352780 $Y=456700
X3138 1969 2 1957 1972 1 NR2 $T=354020 467160 0 0 $X=354020 $Y=466780
X3139 1973 2 1953 1980 1 NR2 $T=354020 487320 1 0 $X=354020 $Y=481900
X3140 1969 2 1968 1980 1 NR2 $T=354020 487320 0 0 $X=354020 $Y=486940
X3141 1803 2 147 1989 1 NR2 $T=355260 376440 0 0 $X=355260 $Y=376060
X3142 107 2 149 117 1 NR2 $T=355880 366360 0 0 $X=355880 $Y=365980
X3143 1969 2 1928 1995 1 NR2 $T=355880 457080 0 0 $X=355880 $Y=456700
X3144 1967 2 2017 2015 1 NR2 $T=357740 436920 1 0 $X=357740 $Y=431500
X3145 1969 2 1981 2015 1 NR2 $T=357740 457080 1 0 $X=357740 $Y=451660
X3146 2023 2 2007 1972 1 NR2 $T=360220 467160 1 180 $X=358360 $Y=466780
X3147 1967 2 2018 1995 1 NR2 $T=359600 447000 1 0 $X=359600 $Y=441580
X3148 2023 2 1946 2015 1 NR2 $T=360840 457080 1 0 $X=360840 $Y=451660
X3149 1973 2 2022 2032 1 NR2 $T=361460 477240 1 0 $X=361460 $Y=471820
X3150 2034 2 2016 156 1 NR2 $T=364560 386520 0 180 $X=362700 $Y=381100
X3151 1972 2 2009 2045 1 NR2 $T=363320 447000 0 0 $X=363320 $Y=446620
X3152 2023 2 2066 1995 1 NR2 $T=366420 477240 0 180 $X=364560 $Y=471820
X3153 1969 2 2038 2032 1 NR2 $T=365180 487320 0 0 $X=365180 $Y=486940
X3154 2015 2 2058 2045 1 NR2 $T=366420 436920 1 0 $X=366420 $Y=431500
X3155 2061 2 2030 2037 1 NR2 $T=368280 447000 1 180 $X=366420 $Y=446620
X3156 1972 2 2072 2037 1 NR2 $T=368900 447000 0 0 $X=368900 $Y=446620
X3157 1967 2 2079 2096 1 NR2 $T=370140 436920 1 0 $X=370140 $Y=431500
X3158 2092 2 1964 2062 1 NR2 $T=372000 487320 0 180 $X=370140 $Y=481900
X3159 1973 2 2077 2098 1 NR2 $T=370760 477240 0 0 $X=370760 $Y=476860
X3160 2106 2 2086 2045 1 NR2 $T=375100 457080 1 180 $X=373240 $Y=456700
X3161 2046 2 2094 2096 1 NR2 $T=373860 436920 0 0 $X=373860 $Y=436540
X3162 2023 2 2109 2098 1 NR2 $T=375720 487320 0 180 $X=373860 $Y=481900
X3163 2119 2 2060 2045 1 NR2 $T=376960 457080 1 180 $X=375100 $Y=456700
X3164 2119 2 1993 2128 1 NR2 $T=375720 457080 1 0 $X=375720 $Y=451660
X3165 2130 2 2057 2015 1 NR2 $T=377580 467160 1 180 $X=375720 $Y=466780
X3166 2023 2 2122 1980 1 NR2 $T=375720 487320 1 0 $X=375720 $Y=481900
X3167 2106 2 2136 2037 1 NR2 $T=377580 457080 0 0 $X=377580 $Y=456700
X3168 2061 2 2156 2045 1 NR2 $T=381300 457080 0 180 $X=379440 $Y=451660
X3169 2130 2 2142 2062 1 NR2 $T=379440 487320 1 0 $X=379440 $Y=481900
X3170 2119 2 2140 2149 1 NR2 $T=382540 426840 0 180 $X=380680 $Y=421420
X3171 2061 2 2162 2128 1 NR2 $T=380680 436920 0 0 $X=380680 $Y=436540
X3172 2092 2 2150 2015 1 NR2 $T=380680 467160 0 0 $X=380680 $Y=466780
X3173 2092 2 2164 1980 1 NR2 $T=380680 487320 0 0 $X=380680 $Y=486940
X3174 2106 2 2146 2149 1 NR2 $T=381300 426840 0 0 $X=381300 $Y=426460
X3175 2061 2 2129 2153 1 NR2 $T=382540 436920 1 0 $X=382540 $Y=431500
X3176 2119 2 2158 2037 1 NR2 $T=384400 457080 0 180 $X=382540 $Y=451660
X3177 2130 2 2159 2184 1 NR2 $T=382540 487320 1 0 $X=382540 $Y=481900
X3178 2181 2 2097 2128 1 NR2 $T=386260 426840 1 180 $X=384400 $Y=426460
X3179 2119 2 2205 2153 1 NR2 $T=384400 436920 0 0 $X=384400 $Y=436540
X3180 2130 2 2188 2182 1 NR2 $T=384400 467160 0 0 $X=384400 $Y=466780
X3181 2092 2 2088 2184 1 NR2 $T=384400 497400 1 0 $X=384400 $Y=491980
X3182 2171 2 2202 2165 1 NR2 $T=384400 507480 0 0 $X=384400 $Y=507100
X3183 174 2 2127 2186 1 NR2 $T=388120 436920 0 180 $X=386260 $Y=431500
X3184 2182 2 2183 2062 1 NR2 $T=386260 477240 0 0 $X=386260 $Y=476860
X3185 2182 2 2069 2194 1 NR2 $T=386260 487320 0 0 $X=386260 $Y=486940
X3186 2190 2 2175 2198 1 NR2 $T=387500 406680 0 0 $X=387500 $Y=406300
X3187 2181 2 2179 176 1 NR2 $T=388120 396600 1 0 $X=388120 $Y=391180
X3188 2198 2 2180 176 1 NR2 $T=388120 416760 1 0 $X=388120 $Y=411340
X3189 2194 2 2208 2062 1 NR2 $T=389980 487320 1 180 $X=388120 $Y=486940
X3190 2091 2 2193 2216 1 NR2 $T=389360 436920 1 0 $X=389360 $Y=431500
X3191 2190 2 2215 2222 1 NR2 $T=389980 406680 1 0 $X=389980 $Y=401260
X3192 2130 2 2206 2061 1 NR2 $T=389980 467160 1 0 $X=389980 $Y=461740
X3193 178 2 2210 2145 1 NR2 $T=390600 386520 0 0 $X=390600 $Y=386140
X3194 179 2 2204 182 1 NR2 $T=391220 386520 1 0 $X=391220 $Y=381100
X3195 2181 2 2191 183 1 NR2 $T=391220 396600 1 0 $X=391220 $Y=391180
X3196 2225 2 2192 178 1 NR2 $T=393080 396600 1 180 $X=391220 $Y=396220
X3197 174 2 2207 2145 1 NR2 $T=394320 386520 1 180 $X=392460 $Y=386140
X3198 2181 2 2230 2153 1 NR2 $T=393080 416760 1 0 $X=393080 $Y=411340
X3199 2216 2 2217 2186 1 NR2 $T=394940 436920 1 180 $X=393080 $Y=436540
X3200 2046 2 2242 2091 1 NR2 $T=395560 436920 0 180 $X=393700 $Y=431500
X3201 2216 2 2248 2187 1 NR2 $T=393700 457080 1 0 $X=393700 $Y=451660
X3202 2246 2 2235 2202 1 NR2 $T=395560 507480 1 180 $X=393700 $Y=507100
X3203 2092 2 2238 2032 1 NR2 $T=394320 487320 0 0 $X=394320 $Y=486940
X3204 187 2 2244 174 1 NR2 $T=396800 386520 1 180 $X=394940 $Y=386140
X3205 2236 2 2241 2153 1 NR2 $T=396800 416760 0 180 $X=394940 $Y=411340
X3206 2198 2 2247 2251 1 NR2 $T=395560 406680 1 0 $X=395560 $Y=401260
X3207 2046 2 2237 2186 1 NR2 $T=397420 426840 0 180 $X=395560 $Y=421420
X3208 2182 2 2255 2187 1 NR2 $T=396180 457080 0 0 $X=396180 $Y=456700
X3209 185 2 2259 2145 1 NR2 $T=396800 386520 0 0 $X=396800 $Y=386140
X3210 2046 2 2253 185 1 NR2 $T=396800 416760 0 0 $X=396800 $Y=416380
X3211 2225 2 2275 2216 1 NR2 $T=398660 436920 0 180 $X=396800 $Y=431500
X3212 2119 2 2231 2251 1 NR2 $T=397420 426840 1 0 $X=397420 $Y=421420
X3213 2184 2 2264 1980 1 NR2 $T=400520 487320 1 180 $X=398660 $Y=486940
X3214 2257 2 2246 2229 1 NR2 $T=398660 517560 1 0 $X=398660 $Y=512140
X3215 196 2 2274 182 1 NR2 $T=401140 386520 1 180 $X=399280 $Y=386140
X3216 2198 2 2287 2149 1 NR2 $T=399280 426840 0 0 $X=399280 $Y=426460
X3217 2236 2 2277 2222 1 NR2 $T=401140 447000 1 180 $X=399280 $Y=446620
X3218 196 2 2272 2145 1 NR2 $T=401760 416760 1 180 $X=399900 $Y=416380
X3219 2282 2 2232 2251 1 NR2 $T=402380 426840 0 180 $X=400520 $Y=421420
X3220 1967 2 2276 2236 1 NR2 $T=400520 447000 1 0 $X=400520 $Y=441580
X3221 196 2 2281 2288 1 NR2 $T=401140 386520 1 0 $X=401140 $Y=381100
X3222 2245 2 2301 2260 1 NR2 $T=403620 436920 1 180 $X=401760 $Y=436540
X3223 2245 2 2293 2222 1 NR2 $T=404240 447000 1 180 $X=402380 $Y=446620
X3224 174 2 2273 186 1 NR2 $T=403000 376440 1 0 $X=403000 $Y=371020
X3225 2298 2 2286 183 1 NR2 $T=404860 376440 0 0 $X=404860 $Y=376060
X3226 205 2 2262 2251 1 NR2 $T=407340 366360 1 180 $X=405480 $Y=365980
X3227 2267 2 2324 2128 1 NR2 $T=407340 447000 1 180 $X=405480 $Y=446620
X3228 2267 2 2310 2292 1 NR2 $T=405480 467160 1 0 $X=405480 $Y=461740
X3229 2292 2 2306 2149 1 NR2 $T=407960 426840 0 180 $X=406100 $Y=421420
X3230 2317 2 2296 2128 1 NR2 $T=407960 436920 1 180 $X=406100 $Y=436540
X3231 2181 2 2326 2251 1 NR2 $T=409200 396600 0 180 $X=407340 $Y=391180
X3232 2198 2 2341 183 1 NR2 $T=407340 396600 0 0 $X=407340 $Y=396220
X3233 2236 2 2328 2187 1 NR2 $T=407340 457080 1 0 $X=407340 $Y=451660
X3234 206 2 207 2298 1 NR2 $T=409820 366360 1 180 $X=407960 $Y=365980
X3235 205 2 2321 2288 1 NR2 $T=409820 376440 0 180 $X=407960 $Y=371020
X3236 2317 2 2320 197 1 NR2 $T=407960 477240 1 0 $X=407960 $Y=471820
X3237 2298 2 2325 176 1 NR2 $T=409200 376440 0 0 $X=409200 $Y=376060
X3238 196 2 2355 171 1 NR2 $T=409200 386520 1 0 $X=409200 $Y=381100
X3239 2267 2 2327 186 1 NR2 $T=411060 426840 0 180 $X=409200 $Y=421420
X3240 2298 2 2315 171 1 NR2 $T=409820 406680 0 0 $X=409820 $Y=406300
X3241 2267 2 2335 171 1 NR2 $T=410440 406680 1 0 $X=410440 $Y=401260
X3242 2282 2 2336 176 1 NR2 $T=410440 416760 1 0 $X=410440 $Y=411340
X3243 2190 2 2340 2181 1 NR2 $T=412920 396600 0 180 $X=411060 $Y=391180
X3244 2317 2 2345 2292 1 NR2 $T=412920 457080 0 180 $X=411060 $Y=451660
X3245 2194 2 2351 188 1 NR2 $T=411060 487320 0 0 $X=411060 $Y=486940
X3246 2222 2 2361 176 1 NR2 $T=412920 396600 0 0 $X=412920 $Y=396220
X3247 206 2 2348 2282 1 NR2 $T=414780 406680 1 180 $X=412920 $Y=406300
X3248 183 2 2349 2282 1 NR2 $T=414780 426840 0 180 $X=412920 $Y=421420
X3249 183 2 2350 2222 1 NR2 $T=414780 426840 1 180 $X=412920 $Y=426460
X3250 2194 2 2330 197 1 NR2 $T=414780 477240 0 180 $X=412920 $Y=471820
X3251 2194 2 2366 210 1 NR2 $T=414780 487320 0 0 $X=414780 $Y=486940
X3252 2184 2 2363 210 1 NR2 $T=414780 497400 0 0 $X=414780 $Y=497020
X3253 2317 2 2365 188 1 NR2 $T=416020 477240 1 0 $X=416020 $Y=471820
X3254 2184 2 2377 188 1 NR2 $T=416640 487320 1 0 $X=416640 $Y=481900
X3255 2317 2 2383 2282 1 NR2 $T=417880 477240 0 0 $X=417880 $Y=476860
X3256 107 2 2405 217 1 NR2 $T=422840 366360 0 0 $X=422840 $Y=365980
X3257 2402 2 2034 2413 1 NR2 $T=424700 396600 0 0 $X=424700 $Y=396220
X3258 2399 2 2413 2421 1 NR2 $T=429040 406680 0 180 $X=427180 $Y=401260
X3259 228 2 2427 2415 1 NR2 $T=429040 436920 0 0 $X=429040 $Y=436540
X3260 2421 2 2466 233 1 NR2 $T=432140 406680 0 0 $X=432140 $Y=406300
X3261 2435 2 2450 2458 1 NR2 $T=432140 527640 0 0 $X=432140 $Y=527260
X3262 2464 2 2438 2452 1 NR2 $T=435240 426840 0 180 $X=433380 $Y=421420
X3263 2420 2 2448 233 1 NR2 $T=434000 376440 0 0 $X=434000 $Y=376060
X3264 240 2 2497 233 1 NR2 $T=437720 386520 0 0 $X=437720 $Y=386140
X3265 246 2 2503 2415 1 NR2 $T=442060 447000 0 180 $X=440200 $Y=441580
X3266 2533 2 2512 233 1 NR2 $T=445160 386520 1 180 $X=443300 $Y=386140
X3267 2556 2 2515 2518 1 NR2 $T=445780 436920 0 180 $X=443920 $Y=431500
X3268 2530 2 2479 2518 1 NR2 $T=446400 426840 0 180 $X=444540 $Y=421420
X3269 2519 2 2500 2547 1 NR2 $T=444540 457080 0 0 $X=444540 $Y=456700
X3270 2536 2 2457 255 1 NR2 $T=445780 487320 0 0 $X=445780 $Y=486940
X3271 2555 2 2563 2547 1 NR2 $T=448260 467160 1 0 $X=448260 $Y=461740
X3272 2563 2 2571 2542 1 NR2 $T=451980 447000 1 180 $X=450120 $Y=446620
X3273 2557 2 255 193 1 NR2 $T=451980 487320 1 0 $X=451980 $Y=481900
X3274 2575 2 2601 2594 1 NR2 $T=455080 457080 1 0 $X=455080 $Y=451660
X3275 2541 2 2615 2609 1 NR2 $T=456940 416760 0 0 $X=456940 $Y=416380
X3276 2611 2 2386 2605 1 NR2 $T=459420 497400 0 180 $X=457560 $Y=491980
X3277 2595 2 2596 2620 1 NR2 $T=458800 487320 1 0 $X=458800 $Y=481900
X3278 2519 2 2608 268 1 NR2 $T=460040 467160 0 0 $X=460040 $Y=466780
X3279 2625 2 2628 2610 1 NR2 $T=462520 447000 0 180 $X=460660 $Y=441580
X3280 2555 2 2662 268 1 NR2 $T=460660 467160 1 0 $X=460660 $Y=461740
X3281 2630 2 2584 2562 1 NR2 $T=463140 487320 1 180 $X=461280 $Y=486940
X3282 2637 2 2644 271 1 NR2 $T=462520 527640 1 0 $X=462520 $Y=522220
X3283 2670 2 2595 2586 1 NR2 $T=468100 477240 1 180 $X=466240 $Y=476860
X3284 2645 2 2667 2604 1 NR2 $T=466240 487320 1 0 $X=466240 $Y=481900
X3285 276 2 2671 282 1 NR2 $T=467480 517560 1 0 $X=467480 $Y=512140
X3286 2617 2 2670 281 1 NR2 $T=468100 477240 0 0 $X=468100 $Y=476860
X3287 2659 2 2635 282 1 NR2 $T=468100 517560 0 0 $X=468100 $Y=517180
X3288 278 2 2651 279 1 NR2 $T=468100 527640 1 0 $X=468100 $Y=522220
X3289 286 2 2668 2659 1 NR2 $T=469960 517560 1 0 $X=469960 $Y=512140
X3290 2547 2 2679 268 1 NR2 $T=472440 467160 0 180 $X=470580 $Y=461740
X3291 2659 2 2691 2637 1 NR2 $T=471820 517560 0 0 $X=471820 $Y=517180
X3292 2642 2 2693 2702 1 NR2 $T=472440 396600 0 0 $X=472440 $Y=396220
X3293 2698 2 281 2707 1 NR2 $T=473060 487320 0 0 $X=473060 $Y=486940
X3294 286 2 2696 271 1 NR2 $T=474300 527640 0 0 $X=474300 $Y=527260
X3295 278 2 2715 2637 1 NR2 $T=474920 517560 0 0 $X=474920 $Y=517180
X3296 2698 2 2721 2605 1 NR2 $T=475540 487320 0 0 $X=475540 $Y=486940
X3297 2519 2 2717 279 1 NR2 $T=476780 477240 0 0 $X=476780 $Y=476860
X3298 286 2 2733 278 1 NR2 $T=476780 527640 1 0 $X=476780 $Y=522220
X3299 278 2 2725 282 1 NR2 $T=478640 527640 1 180 $X=476780 $Y=527260
X3300 279 2 2710 2742 1 NR2 $T=478640 487320 1 0 $X=478640 $Y=481900
X3301 258 2 2748 2684 1 NR2 $T=482360 487320 0 180 $X=480500 $Y=481900
X3302 276 2 2751 2637 1 NR2 $T=480500 517560 0 0 $X=480500 $Y=517180
X3303 276 2 2738 279 1 NR2 $T=482360 527640 0 180 $X=480500 $Y=522220
X3304 2742 2 2761 278 1 NR2 $T=483600 507480 1 180 $X=481740 $Y=507100
X3305 2731 2 2771 2561 1 NR2 $T=482360 487320 1 0 $X=482360 $Y=481900
X3306 2637 2 298 300 1 NR2 $T=482360 537720 1 0 $X=482360 $Y=532300
X3307 2697 2 2757 2772 1 NR2 $T=482980 376440 1 0 $X=482980 $Y=371020
X3308 2778 2 2743 302 1 NR2 $T=486080 537720 0 180 $X=484220 $Y=532300
X3309 297 2 2776 2760 1 NR2 $T=486080 487320 0 0 $X=486080 $Y=486940
X3310 306 2 310 311 1 NR2 $T=487320 366360 0 0 $X=487320 $Y=365980
X3311 2742 2 2791 2659 1 NR2 $T=489180 517560 0 180 $X=487320 $Y=512140
X3312 2729 2 2799 2802 1 NR2 $T=489180 416760 1 0 $X=489180 $Y=411340
X3313 2742 2 2794 2760 1 NR2 $T=489180 487320 0 0 $X=489180 $Y=486940
X3314 2778 2 2758 2795 1 NR2 $T=491040 497400 1 180 $X=489180 $Y=497020
X3315 2778 2 2777 317 1 NR2 $T=491040 527640 0 0 $X=491040 $Y=527260
X3316 2810 2 2812 2817 1 NR2 $T=491660 436920 0 0 $X=491660 $Y=436540
X3317 2778 2 2832 304 1 NR2 $T=492900 527640 1 0 $X=492900 $Y=522220
X3318 2844 2 2849 2705 1 NR2 $T=496620 416760 0 0 $X=496620 $Y=416380
X3319 2705 2 2892 2907 1 NR2 $T=504680 406680 0 0 $X=504680 $Y=406300
X3320 2919 2 2826 2871 1 NR2 $T=508400 497400 1 180 $X=506540 $Y=497020
X3321 2932 2 2885 2852 1 NR2 $T=509020 497400 0 180 $X=507160 $Y=491980
X3322 2921 2 2851 2871 1 NR2 $T=508400 497400 0 0 $X=508400 $Y=497020
X3323 2937 2 2934 2852 1 NR2 $T=510260 507480 0 180 $X=508400 $Y=502060
X3324 2921 2 2911 2852 1 NR2 $T=508400 507480 0 0 $X=508400 $Y=507100
X3325 2919 2 2928 2852 1 NR2 $T=508400 517560 1 0 $X=508400 $Y=512140
X3326 2930 2 2929 2944 1 NR2 $T=509020 376440 1 0 $X=509020 $Y=371020
X3327 2763 2 2935 2880 1 NR2 $T=509020 416760 0 0 $X=509020 $Y=416380
X3328 2932 2 2838 2871 1 NR2 $T=512120 497400 0 180 $X=510260 $Y=491980
X3329 2870 2 2988 2802 1 NR2 $T=510880 406680 0 0 $X=510880 $Y=406300
X3330 2937 2 2916 2871 1 NR2 $T=512740 507480 0 180 $X=510880 $Y=502060
X3331 2855 2 341 2753 1 NR2 $T=513980 426840 0 180 $X=512120 $Y=421420
X3332 2919 2 338 2968 1 NR2 $T=512120 517560 0 0 $X=512120 $Y=517180
X3333 2800 2 340 2940 1 NR2 $T=512740 406680 1 0 $X=512740 $Y=401260
X3334 2901 2 2993 2920 1 NR2 $T=513980 416760 1 0 $X=513980 $Y=411340
X3335 2853 2 2983 2919 1 NR2 $T=515840 517560 1 180 $X=513980 $Y=517180
X3336 3001 2 2986 2920 1 NR2 $T=517080 406680 0 180 $X=515220 $Y=401260
X3337 2940 2 2930 3013 1 NR2 $T=515840 376440 1 0 $X=515840 $Y=371020
X3338 2954 2 3002 2920 1 NR2 $T=517700 416760 0 180 $X=515840 $Y=411340
X3339 2937 2 348 2968 1 NR2 $T=515840 507480 0 0 $X=515840 $Y=507100
X3340 2802 2 3008 2940 1 NR2 $T=517080 406680 1 0 $X=517080 $Y=401260
X3341 2853 2 357 2921 1 NR2 $T=518940 517560 0 0 $X=518940 $Y=517180
X3342 2853 2 356 2932 1 NR2 $T=519560 507480 0 0 $X=519560 $Y=507100
X3343 2940 2 3037 3036 1 NR2 $T=520180 396600 0 0 $X=520180 $Y=396220
X3344 2921 2 2909 2968 1 NR2 $T=520180 517560 1 0 $X=520180 $Y=512140
X3345 2932 2 3046 2968 1 NR2 $T=523280 507480 1 180 $X=521420 $Y=507100
X3346 2940 2 3058 3059 1 NR2 $T=522660 376440 1 0 $X=522660 $Y=371020
X3347 2940 2 3052 3071 1 NR2 $T=522660 396600 1 0 $X=522660 $Y=391180
X3348 3037 2 3072 3083 1 NR2 $T=524520 416760 1 0 $X=524520 $Y=411340
X3349 2729 2 3081 3093 1 NR2 $T=525140 497400 0 0 $X=525140 $Y=497020
X3350 3110 2 3140 3052 1 NR2 $T=530100 396600 1 0 $X=530100 $Y=391180
X3351 3117 2 3150 3137 1 NR2 $T=535060 497400 1 180 $X=533200 $Y=497020
X3352 3159 2 3142 3119 1 NR2 $T=535680 497400 0 180 $X=533820 $Y=491980
X3353 3220 2 3202 3203 1 NR2 $T=542500 447000 0 180 $X=540640 $Y=441580
X3354 3234 2 3230 3195 1 NR2 $T=545600 436920 1 180 $X=543740 $Y=436540
X3355 399 2 393 3257 1 NR2 $T=551800 396600 0 180 $X=549940 $Y=391180
X3356 385 2 3258 3275 1 NR2 $T=550560 376440 1 0 $X=550560 $Y=371020
X3357 3310 2 3262 3285 1 NR2 $T=555520 487320 0 180 $X=553660 $Y=481900
X3358 3314 2 3301 3305 1 NR2 $T=558000 467160 1 180 $X=556140 $Y=466780
X3359 3310 2 3290 3314 1 NR2 $T=556760 487320 1 0 $X=556760 $Y=481900
X3360 3338 2 3274 3329 1 NR2 $T=562340 467160 1 180 $X=560480 $Y=466780
X3361 3342 2 3326 3348 1 NR2 $T=562340 426840 1 0 $X=562340 $Y=421420
X3362 3328 2 3352 3325 1 NR2 $T=562340 447000 1 0 $X=562340 $Y=441580
X3363 3309 2 3357 3349 1 NR2 $T=565440 467160 0 180 $X=563580 $Y=461740
X3364 3314 2 3367 3329 1 NR2 $T=563580 467160 0 0 $X=563580 $Y=466780
X3365 3317 2 3358 3329 1 NR2 $T=564820 477240 0 0 $X=564820 $Y=476860
X3366 3310 2 3355 3329 1 NR2 $T=565440 487320 0 0 $X=565440 $Y=486940
X3367 3372 2 3371 3317 1 NR2 $T=568540 477240 1 180 $X=566680 $Y=476860
X3368 3374 2 3379 3351 1 NR2 $T=569160 436920 1 180 $X=567300 $Y=436540
X3369 3372 2 3378 3305 1 NR2 $T=567920 487320 1 0 $X=567920 $Y=481900
X3370 3369 2 3340 3384 1 NR2 $T=569160 416760 0 0 $X=569160 $Y=416380
X3371 3373 2 3386 3349 1 NR2 $T=570400 497400 0 0 $X=570400 $Y=497020
X3372 3310 2 3411 3349 1 NR2 $T=571640 507480 0 0 $X=571640 $Y=507100
X3373 433 2 3416 424 1 NR2 $T=575980 527640 1 180 $X=574120 $Y=527260
X3374 426 2 3426 429 1 NR2 $T=575980 366360 0 0 $X=575980 $Y=365980
X3375 3428 2 3420 2421 1 NR2 $T=577840 416760 1 180 $X=575980 $Y=416380
X3376 3428 2 3421 2530 1 NR2 $T=577840 426840 0 180 $X=575980 $Y=421420
X3377 3309 2 3432 3429 1 NR2 $T=575980 467160 1 0 $X=575980 $Y=461740
X3378 3338 2 3350 3429 1 NR2 $T=575980 467160 0 0 $X=575980 $Y=466780
X3379 3338 2 3425 430 1 NR2 $T=576600 477240 0 0 $X=576600 $Y=476860
X3380 3317 2 3423 430 1 NR2 $T=576600 487320 0 0 $X=576600 $Y=486940
X3381 3317 2 3440 3408 1 NR2 $T=577840 487320 1 0 $X=577840 $Y=481900
X3382 3317 2 3448 3429 1 NR2 $T=578460 477240 1 0 $X=578460 $Y=471820
X3383 3428 2 3443 3115 1 NR2 $T=581560 416760 0 180 $X=579700 $Y=411340
X3384 440 2 439 213 1 NR2 $T=582800 366360 1 180 $X=580940 $Y=365980
X3385 3305 2 3434 3429 1 NR2 $T=581560 487320 1 0 $X=581560 $Y=481900
X3386 437 2 3467 430 1 NR2 $T=581560 487320 0 0 $X=581560 $Y=486940
X3387 3159 2 3401 444 1 NR2 $T=581560 497400 1 0 $X=581560 $Y=491980
X3388 3441 2 3459 442 1 NR2 $T=584660 366360 1 180 $X=582800 $Y=365980
X3389 3441 2 3454 323 1 NR2 $T=585280 376440 0 180 $X=583420 $Y=371020
X3390 3441 2 3463 2420 1 NR2 $T=585280 386520 1 180 $X=583420 $Y=386140
X3391 3441 2 3464 2533 1 NR2 $T=585280 406680 0 180 $X=583420 $Y=401260
X3392 3441 2 3493 240 1 NR2 $T=585280 406680 1 180 $X=583420 $Y=406300
X3393 3159 2 3480 453 1 NR2 $T=584040 497400 0 0 $X=584040 $Y=497020
X3394 3453 2 3460 3450 1 NR2 $T=587140 447000 1 180 $X=585280 $Y=446620
X3395 3309 2 3490 430 1 NR2 $T=587760 487320 1 0 $X=587760 $Y=481900
X3396 3314 2 3494 3429 1 NR2 $T=589000 467160 0 0 $X=589000 $Y=466780
X3397 3519 2 3495 3505 1 NR2 $T=592100 406680 0 180 $X=590240 $Y=401260
X3398 3485 2 3502 3456 1 NR2 $T=590240 447000 1 0 $X=590240 $Y=441580
X3399 3418 2 3403 3429 1 NR2 $T=592100 507480 1 180 $X=590240 $Y=507100
X3400 449 2 3499 444 1 NR2 $T=590240 537720 1 0 $X=590240 $Y=532300
X3401 3338 2 3543 3557 1 NR2 $T=593960 467160 0 0 $X=593960 $Y=466780
X3402 3563 2 3521 3549 1 NR2 $T=598920 406680 1 180 $X=597060 $Y=406300
X3403 3373 2 3564 3305 1 NR2 $T=599540 477240 0 180 $X=597680 $Y=471820
X3404 3562 2 3561 3458 1 NR2 $T=599540 507480 1 180 $X=597680 $Y=507100
X3405 3428 2 3570 2556 1 NR2 $T=601400 436920 1 180 $X=599540 $Y=436540
X3406 3572 2 3594 3408 1 NR2 $T=602640 497400 0 0 $X=602640 $Y=497020
X3407 3593 2 3563 3583 1 NR2 $T=605120 406680 0 180 $X=603260 $Y=401260
X3408 450 2 3616 3614 1 NR2 $T=604500 497400 1 0 $X=604500 $Y=491980
X3409 3586 2 3602 3574 1 NR2 $T=605120 507480 0 0 $X=605120 $Y=507100
X3410 3620 2 3578 3598 1 NR2 $T=608220 447000 0 180 $X=606360 $Y=441580
X3411 463 2 3615 3614 1 NR2 $T=608840 487320 1 180 $X=606980 $Y=486940
X3412 3590 2 3629 3636 1 NR2 $T=608220 457080 1 0 $X=608220 $Y=451660
X3413 3658 2 3605 3590 1 NR2 $T=610080 457080 1 180 $X=608220 $Y=456700
X3414 450 2 3622 3630 1 NR2 $T=608220 477240 1 0 $X=608220 $Y=471820
X3415 403 2 3624 423 1 NR2 $T=608220 527640 1 0 $X=608220 $Y=522220
X3416 3373 2 3643 465 1 NR2 $T=610080 507480 1 0 $X=610080 $Y=502060
X3417 3617 2 3632 444 1 NR2 $T=610080 527640 0 0 $X=610080 $Y=527260
X3418 463 2 3648 430 1 NR2 $T=613800 527640 1 180 $X=611940 $Y=527260
X3419 3557 2 3653 3630 1 NR2 $T=614420 477240 0 180 $X=612560 $Y=471820
X3420 444 2 3677 3659 1 NR2 $T=613180 517560 1 0 $X=613180 $Y=512140
X3421 3557 2 3685 3590 1 NR2 $T=613800 467160 0 0 $X=613800 $Y=466780
X3422 453 2 3663 3659 1 NR2 $T=615660 527640 1 180 $X=613800 $Y=527260
X3423 3666 2 3689 3590 1 NR2 $T=614420 477240 1 0 $X=614420 $Y=471820
X3424 3671 2 3541 3657 1 NR2 $T=615040 436920 1 0 $X=615040 $Y=431500
X3425 3630 2 3682 3659 1 NR2 $T=615040 487320 0 0 $X=615040 $Y=486940
X3426 3658 2 3688 3630 1 NR2 $T=617520 467160 0 180 $X=615660 $Y=461740
X3427 463 2 3691 3658 1 NR2 $T=615660 497400 1 0 $X=615660 $Y=491980
X3428 453 2 3702 450 1 NR2 $T=618140 497400 1 180 $X=616280 $Y=497020
X3429 3590 2 3704 3659 1 NR2 $T=617520 487320 0 0 $X=617520 $Y=486940
X3430 3658 2 3700 3614 1 NR2 $T=618140 467160 0 0 $X=618140 $Y=466780
X3431 3692 2 3671 3723 1 NR2 $T=622480 436920 1 0 $X=622480 $Y=431500
X3432 3745 2 3526 3731 1 NR2 $T=626200 426840 0 0 $X=626200 $Y=426460
X3433 3737 2 3748 3718 1 NR2 $T=626200 447000 1 0 $X=626200 $Y=441580
X3434 3716 2 3755 3699 1 NR2 $T=627440 447000 0 0 $X=627440 $Y=446620
X3435 3793 2 3657 3772 1 NR2 $T=634880 436920 1 180 $X=633020 $Y=436540
X3436 3610 2 3799 480 1 NR2 $T=636120 517560 1 180 $X=634260 $Y=517180
X3437 3788 2 3794 3805 1 NR2 $T=634880 527640 1 0 $X=634880 $Y=522220
X3438 3840 2 3837 3828 1 NR2 $T=643560 447000 1 180 $X=641700 $Y=446620
X3439 3835 2 3850 3817 1 NR2 $T=645420 457080 1 0 $X=645420 $Y=451660
X3440 501 2 3870 3766 1 NR2 $T=647280 517560 1 0 $X=647280 $Y=512140
X3441 499 2 3878 496 1 NR2 $T=647280 537720 1 0 $X=647280 $Y=532300
X3442 3883 2 3886 3871 1 NR2 $T=651000 497400 1 0 $X=651000 $Y=491980
X3443 3847 2 3898 3852 1 NR2 $T=654100 477240 1 180 $X=652240 $Y=476860
X3444 3902 2 3913 3904 1 NR2 $T=656580 527640 0 180 $X=654720 $Y=522220
X3445 3912 2 3906 3890 1 NR2 $T=657820 487320 1 0 $X=657820 $Y=481900
X3446 602 2 4219 598 1 NR2 $T=737800 426840 1 180 $X=735940 $Y=426460
X3447 602 2 4336 605 1 NR2 $T=737800 426840 1 0 $X=737800 $Y=421420
X3448 602 2 4354 609 1 NR2 $T=742760 457080 0 0 $X=742760 $Y=456700
X3449 4353 2 4363 609 1 NR2 $T=746480 517560 0 180 $X=744620 $Y=512140
X3450 616 2 4365 609 1 NR2 $T=747100 457080 1 180 $X=745240 $Y=456700
X3451 619 2 4371 609 1 NR2 $T=748340 507480 0 180 $X=746480 $Y=502060
X3452 4390 2 4372 598 1 NR2 $T=750200 477240 1 180 $X=748340 $Y=476860
X3453 619 2 4380 598 1 NR2 $T=748960 467160 0 0 $X=748960 $Y=466780
X3454 619 2 4389 605 1 NR2 $T=748960 487320 0 0 $X=748960 $Y=486940
X3455 4353 2 4387 598 1 NR2 $T=750820 537720 0 180 $X=748960 $Y=532300
X3456 624 2 4392 598 1 NR2 $T=752680 426840 0 180 $X=750820 $Y=421420
X3457 4388 2 4402 598 1 NR2 $T=753920 416760 1 180 $X=752060 $Y=416380
X3458 619 2 4746 701 1 NR2 $T=827700 467160 0 0 $X=827700 $Y=466780
X3459 4353 2 4755 701 1 NR2 $T=830180 507480 1 0 $X=830180 $Y=502060
X3460 4388 2 4762 701 1 NR2 $T=832040 436920 1 0 $X=832040 $Y=431500
X3461 602 2 4774 701 1 NR2 $T=837620 436920 0 180 $X=835760 $Y=431500
X3462 602 2 4916 765 1 NR2 $T=859940 436920 0 0 $X=859940 $Y=436540
X3463 4940 2 4947 766 1 NR2 $T=866140 426840 0 0 $X=866140 $Y=426460
X3464 4390 2 5007 803 1 NR2 $T=880400 477240 0 0 $X=880400 $Y=476860
X3465 4895 2 5057 803 1 NR2 $T=889080 477240 1 0 $X=889080 $Y=471820
X3466 4940 2 5054 803 1 NR2 $T=890320 426840 0 0 $X=890320 $Y=426460
X3467 624 2 5069 803 1 NR2 $T=894040 426840 1 180 $X=892180 $Y=426460
X3468 4353 2 5449 939 1 NR2 $T=975880 497400 0 0 $X=975880 $Y=497020
X3469 4895 2 5461 939 1 NR2 $T=978980 467160 1 0 $X=978980 $Y=461740
X3470 4388 2 5479 939 1 NR2 $T=981460 416760 0 0 $X=981460 $Y=416380
X3471 4940 2 5455 939 1 NR2 $T=984560 426840 0 180 $X=982700 $Y=421420
X3472 4895 2 5515 969 1 NR2 $T=987660 487320 0 0 $X=987660 $Y=486940
X3473 4895 2 5555 984 1 NR2 $T=995720 467160 1 0 $X=995720 $Y=461740
X3474 624 2 5563 969 1 NR2 $T=998820 416760 0 0 $X=998820 $Y=416380
X3475 4940 2 5574 969 1 NR2 $T=1002540 426840 0 180 $X=1000680 $Y=421420
X3476 624 2 5614 984 1 NR2 $T=1002540 426840 1 0 $X=1002540 $Y=421420
X3477 1923 231 1 2 INV12CK $T=437100 477240 0 180 $X=427180 $Y=471820
X3478 4582 3926 1 2 INV12CK $T=792980 487320 0 180 $X=783060 $Y=481900
X3479 4582 612 1 2 INV12CK $T=794840 507480 0 180 $X=784920 $Y=502060
X3480 663 4582 1 2 INV12CK $T=795460 497400 0 180 $X=785540 $Y=491980
X3481 4582 4560 1 2 INV12CK $T=799180 497400 0 0 $X=799180 $Y=497020
X3482 953 846 1 2 INV12CK $T=982700 376440 0 0 $X=982700 $Y=376060
X3483 1096 1039 1 2 INV12CK $T=1081900 497400 0 0 $X=1081900 $Y=497020
X3484 1323 1328 2 1 1347 OR2 $T=243660 426840 1 0 $X=243660 $Y=421420
X3485 1366 1301 2 1 1409 OR2 $T=254200 386520 0 0 $X=254200 $Y=386140
X3486 1355 1390 2 1 1418 OR2 $T=257920 447000 0 0 $X=257920 $Y=446620
X3487 1405 1397 2 1 58 OR2 $T=258540 366360 0 0 $X=258540 $Y=365980
X3488 1408 1431 2 1 1475 OR2 $T=265360 477240 1 0 $X=265360 $Y=471820
X3489 1469 1472 2 1 1508 OR2 $T=274040 477240 0 0 $X=274040 $Y=476860
X3490 1522 76 2 1 1538 OR2 $T=283960 507480 0 0 $X=283960 $Y=507100
X3491 95 96 2 1 97 OR2 $T=300700 366360 0 0 $X=300700 $Y=365980
X3492 1885 1898 2 1 1906 OR2 $T=341620 517560 0 0 $X=341620 $Y=517180
X3493 1840 1990 2 1 1989 OR2 $T=355880 386520 0 0 $X=355880 $Y=386140
X3494 2056 2047 2 1 1998 OR2 $T=367040 507480 1 180 $X=364560 $Y=507100
X3495 2314 2319 2 1 2418 OR2 $T=423460 507480 0 0 $X=423460 $Y=507100
X3496 2359 2395 2 1 2429 OR2 $T=426560 507480 0 0 $X=426560 $Y=507100
X3497 2459 2431 2 1 2473 OR2 $T=434000 517560 1 0 $X=434000 $Y=512140
X3498 2474 236 2 1 2490 OR2 $T=435860 527640 0 0 $X=435860 $Y=527260
X3499 2487 2482 2 1 2476 OR2 $T=438960 426840 1 180 $X=436480 $Y=426460
X3500 2555 2519 2 1 2499 OR2 $T=447020 467160 0 180 $X=444540 $Y=461740
X3501 258 2562 2 1 2536 OR2 $T=450740 487320 1 180 $X=448260 $Y=486940
X3502 2561 2562 2 1 259 OR2 $T=449500 487320 1 0 $X=449500 $Y=481900
X3503 2386 258 2 1 2561 OR2 $T=451360 497400 1 0 $X=451360 $Y=491980
X3504 259 2557 2 1 2485 OR2 $T=451980 467160 0 0 $X=451980 $Y=466780
X3505 2611 2613 2 1 2562 OR2 $T=458800 487320 0 0 $X=458800 $Y=486940
X3506 2617 2611 2 1 2645 OR2 $T=460040 477240 0 0 $X=460040 $Y=476860
X3507 2611 2604 2 1 2650 OR2 $T=462520 497400 1 0 $X=462520 $Y=491980
X3508 2643 2588 2 1 2669 OR2 $T=463760 406680 1 0 $X=463760 $Y=401260
X3509 2650 2630 2 1 2684 OR2 $T=465620 487320 0 0 $X=465620 $Y=486940
X3510 2617 2613 2 1 2605 OR2 $T=465620 497400 1 0 $X=465620 $Y=491980
X3511 2711 2716 2 1 2724 OR2 $T=474920 376440 0 0 $X=474920 $Y=376060
X3512 2836 2800 2 1 2918 OR2 $T=504680 396600 0 0 $X=504680 $Y=396220
X3513 2918 2870 2 1 2901 OR2 $T=507160 416760 0 180 $X=504680 $Y=411340
X3514 2729 2834 2 1 2921 OR2 $T=505920 436920 1 0 $X=505920 $Y=431500
X3515 2895 2800 2 1 2938 OR2 $T=507780 396600 0 0 $X=507780 $Y=396220
X3516 2920 2705 2 1 2940 OR2 $T=508400 406680 0 0 $X=508400 $Y=406300
X3517 2753 2729 2 1 2937 OR2 $T=508400 426840 1 0 $X=508400 $Y=421420
X3518 2834 2855 2 1 2932 OR2 $T=508400 436920 1 0 $X=508400 $Y=431500
X3519 2938 2870 2 1 2954 OR2 $T=510260 396600 0 0 $X=510260 $Y=396220
X3520 2954 2763 2 1 2968 OR2 $T=512120 416760 0 0 $X=512120 $Y=416380
X3521 3168 3180 2 1 3067 OR2 $T=539400 396600 0 180 $X=536920 $Y=391180
X3522 3445 3437 2 1 3410 OR2 $T=580940 386520 0 180 $X=578460 $Y=381100
X3523 441 3426 2 1 3437 OR2 $T=582180 376440 1 180 $X=579700 $Y=376060
X3524 3523 451 2 1 3509 OR2 $T=593340 376440 0 0 $X=593340 $Y=376060
X3525 3565 3560 2 1 3528 OR2 $T=600160 396600 0 180 $X=597680 $Y=391180
X3526 3608 3590 2 1 3542 OR2 $T=605120 457080 1 180 $X=602640 $Y=456700
X3527 3608 3557 2 1 3596 OR2 $T=606980 477240 0 180 $X=604500 $Y=471820
X3528 3244 3408 2 1 3609 OR2 $T=604500 487320 0 0 $X=604500 $Y=486940
X3529 3608 3614 2 1 3604 OR2 $T=608220 457080 0 180 $X=605740 $Y=451660
X3530 3244 3418 2 1 3637 OR2 $T=607600 507480 0 0 $X=607600 $Y=507100
X3531 3244 464 2 1 3628 OR2 $T=607600 527640 0 0 $X=607600 $Y=527260
X3532 3642 3635 2 1 3567 OR2 $T=611320 416760 1 180 $X=608840 $Y=416380
X3533 3244 3373 2 1 3639 OR2 $T=608840 487320 0 0 $X=608840 $Y=486940
X3534 3654 3636 2 1 3620 OR2 $T=613800 457080 0 180 $X=611320 $Y=451660
X3535 3678 3664 2 1 3522 OR2 $T=615660 416760 1 180 $X=613180 $Y=416380
X3536 3654 3658 2 1 3674 OR2 $T=613180 457080 0 0 $X=613180 $Y=456700
X3537 3608 3666 2 1 3732 OR2 $T=618760 467160 1 0 $X=618760 $Y=461740
X3538 3659 3608 2 1 3733 OR2 $T=618760 477240 0 0 $X=618760 $Y=476860
X3539 605 4388 2 1 4231 OR2 $T=750820 426840 0 180 $X=748340 $Y=421420
X3540 765 619 2 1 4822 OR2 $T=860560 477240 0 180 $X=858080 $Y=471820
X3541 765 4353 2 1 4841 OR2 $T=859940 517560 1 0 $X=859940 $Y=512140
X3542 766 4353 2 1 4915 OR2 $T=859940 517560 0 0 $X=859940 $Y=517180
X3543 766 4895 2 1 4926 OR2 $T=861800 477240 1 0 $X=861800 $Y=471820
X3544 765 4388 2 1 4886 OR2 $T=866140 426840 1 180 $X=863660 $Y=426460
X3545 766 4388 2 1 4958 OR2 $T=867380 436920 1 0 $X=867380 $Y=431500
X3546 969 4390 2 1 5467 OR2 $T=991380 507480 1 180 $X=988900 $Y=507100
X3547 981 4895 2 1 5489 OR2 $T=992620 487320 0 180 $X=990140 $Y=481900
X3548 981 624 2 1 5444 OR2 $T=993860 426840 0 180 $X=991380 $Y=421420
X3549 981 4390 2 1 5500 OR2 $T=993240 487320 1 0 $X=993240 $Y=481900
X3550 984 4390 2 1 5527 OR2 $T=997580 477240 0 180 $X=995100 $Y=471820
X3551 981 4940 2 1 5511 OR2 $T=996960 426840 1 0 $X=996960 $Y=421420
X3552 984 4940 2 1 5596 OR2 $T=1002540 426840 0 0 $X=1002540 $Y=426460
X3553 1203 1212 1 2 1216 AN2 $T=220720 426840 1 0 $X=220720 $Y=421420
X3554 1237 1224 1 2 1218 AN2 $T=225060 386520 0 180 $X=222580 $Y=381100
X3555 1231 1227 1 2 1204 AN2 $T=225060 467160 1 180 $X=222580 $Y=466780
X3556 1241 1239 1 2 1232 AN2 $T=226920 477240 1 180 $X=224440 $Y=476860
X3557 1293 1255 1 2 1288 AN2 $T=237460 507480 0 180 $X=234980 $Y=502060
X3558 1395 1382 1 2 1403 AN2 $T=256060 527640 1 0 $X=256060 $Y=522220
X3559 1437 1482 1 2 1495 AN2 $T=274040 386520 1 0 $X=274040 $Y=381100
X3560 1473 1482 1 2 1500 AN2 $T=274040 396600 1 0 $X=274040 $Y=391180
X3561 1460 1482 1 2 1497 AN2 $T=275900 406680 1 0 $X=275900 $Y=401260
X3562 1422 1482 1 2 1501 AN2 $T=275900 416760 1 0 $X=275900 $Y=411340
X3563 1490 1482 1 2 1531 AN2 $T=282720 416760 0 0 $X=282720 $Y=416380
X3564 1521 1534 1 2 1543 AN2 $T=284580 457080 1 0 $X=284580 $Y=451660
X3565 1540 1534 1 2 1551 AN2 $T=286440 447000 0 0 $X=286440 $Y=446620
X3566 1563 1534 1 2 1552 AN2 $T=291400 467160 0 180 $X=288920 $Y=461740
X3567 1529 1534 1 2 1586 AN2 $T=291400 436920 1 0 $X=291400 $Y=431500
X3568 1628 1534 1 2 1616 AN2 $T=301940 477240 0 180 $X=299460 $Y=471820
X3569 1653 1674 1 2 1695 AN2 $T=305660 507480 1 0 $X=305660 $Y=502060
X3570 1708 1674 1 2 1725 AN2 $T=309380 507480 1 0 $X=309380 $Y=502060
X3571 1774 1674 1 2 1798 AN2 $T=319920 517560 1 0 $X=319920 $Y=512140
X3572 1922 1933 1 2 1960 AN2 $T=349060 386520 0 0 $X=349060 $Y=386140
X3573 1893 2003 1 2 1976 AN2 $T=358980 527640 0 180 $X=356500 $Y=522220
X3574 1884 2003 1 2 2027 AN2 $T=358980 527640 1 0 $X=358980 $Y=522220
X3575 1978 2003 1 2 2051 AN2 $T=362700 527640 1 0 $X=362700 $Y=522220
X3576 2031 2003 1 2 2074 AN2 $T=367660 517560 0 0 $X=367660 $Y=517180
X3577 2112 2003 1 2 2124 AN2 $T=374480 517560 0 0 $X=374480 $Y=517180
X3578 2209 203 1 2 2333 AN2 $T=405480 527640 0 0 $X=405480 $Y=527260
X3579 2249 203 1 2 2339 AN2 $T=409200 527640 1 0 $X=409200 $Y=522220
X3580 2487 2482 1 2 2495 AN2 $T=438960 426840 0 0 $X=438960 $Y=426460
X3581 2567 2563 1 2 2560 AN2 $T=451360 457080 1 0 $X=451360 $Y=451660
X3582 2590 2607 1 2 260 AN2 $T=457560 426840 1 0 $X=457560 $Y=421420
X3583 2586 2630 1 2 2620 AN2 $T=463140 487320 0 180 $X=460660 $Y=481900
X3584 2643 2588 1 2 2661 AN2 $T=463760 406680 0 0 $X=463760 $Y=406300
X3585 2711 2716 1 2 2750 AN2 $T=474920 386520 1 0 $X=474920 $Y=381100
X3586 2721 2806 1 2 2865 AN2 $T=497240 467160 0 0 $X=497240 $Y=466780
X3587 2860 2824 1 2 2876 AN2 $T=498480 436920 0 0 $X=498480 $Y=436540
X3588 2721 2835 1 2 2878 AN2 $T=499720 467160 0 0 $X=499720 $Y=466780
X3589 2860 2726 1 2 2893 AN2 $T=500960 457080 1 0 $X=500960 $Y=451660
X3590 2860 2864 1 2 2924 AN2 $T=502820 447000 1 0 $X=502820 $Y=441580
X3591 2860 2784 1 2 2902 AN2 $T=502820 447000 0 0 $X=502820 $Y=446620
X3592 2926 2933 1 2 2942 AN2 $T=508400 527640 1 0 $X=508400 $Y=522220
X3593 2969 2942 1 2 2947 AN2 $T=513980 527640 0 180 $X=511500 $Y=522220
X3594 2947 2958 1 2 2965 AN2 $T=511500 527640 0 0 $X=511500 $Y=527260
X3595 2956 2962 1 2 2976 AN2 $T=512120 497400 1 0 $X=512120 $Y=491980
X3596 2970 2991 1 2 2958 AN2 $T=516460 537720 0 180 $X=513980 $Y=532300
X3597 349 2983 1 2 3000 AN2 $T=518320 517560 1 180 $X=515840 $Y=517180
X3598 3011 3018 1 2 3023 AN2 $T=517080 487320 0 0 $X=517080 $Y=486940
X3599 2995 3019 1 2 3024 AN2 $T=517080 507480 1 0 $X=517080 $Y=502060
X3600 3024 3023 1 2 2956 AN2 $T=518940 497400 0 0 $X=518940 $Y=497020
X3601 3034 3032 1 2 2969 AN2 $T=521420 527640 1 180 $X=518940 $Y=527260
X3602 353 3029 1 2 3034 AN2 $T=518940 537720 1 0 $X=518940 $Y=532300
X3603 3077 3085 1 2 3032 AN2 $T=527000 527640 0 180 $X=524520 $Y=522220
X3604 3181 3169 1 2 3194 AN2 $T=538160 416760 0 0 $X=538160 $Y=416380
X3605 3706 3757 1 2 3730 AN2 $T=630540 426840 1 180 $X=628060 $Y=426460
X3606 3823 3849 1 2 3833 AN2 $T=646040 436920 1 180 $X=643560 $Y=436540
X3607 3917 3897 1 2 3895 AN2 $T=654720 467160 0 180 $X=652240 $Y=461740
X3608 137 2 1882 136 1921 1 NR3 $T=350300 366360 1 180 $X=347200 $Y=365980
X3609 144 2 1914 140 1931 1 NR3 $T=354020 366360 1 180 $X=350920 $Y=365980
X3610 1219 1217 1 1286 2 OR2B1S $T=231880 487320 1 0 $X=231880 $Y=481900
X3611 1268 1348 1 1349 2 OR2B1S $T=252340 447000 1 180 $X=249240 $Y=446620
X3612 1319 1359 1 1387 2 OR2B1S $T=251720 507480 0 0 $X=251720 $Y=507100
X3613 1268 1353 1 1417 2 OR2B1S $T=256680 406680 0 0 $X=256680 $Y=406300
X3614 1268 1413 1 1428 2 OR2B1S $T=259160 386520 0 0 $X=259160 $Y=386140
X3615 51 56 1 1457 2 OR2B1S $T=265360 527640 0 0 $X=265360 $Y=527260
X3616 51 70 1 1493 2 OR2B1S $T=274040 537720 1 0 $X=274040 $Y=532300
X3617 2574 2573 1 2551 2 OR2B1S $T=453220 426840 1 0 $X=453220 $Y=421420
X3618 2574 2576 1 2622 2 OR2B1S $T=467480 396600 0 180 $X=464380 $Y=391180
X3619 284 272 1 2677 2 OR2B1S $T=473680 376440 1 180 $X=470580 $Y=376060
X3620 2972 2963 1 2917 2 OR2B1S $T=514600 507480 1 180 $X=511500 $Y=507100
X3621 2957 2965 1 2972 2 OR2B1S $T=512120 517560 1 0 $X=512120 $Y=512140
X3622 3000 2976 1 2957 2 OR2B1S $T=516460 507480 0 180 $X=513360 $Y=502060
X3623 4332 4197 2 1 4349 4351 4123 4216 4320 4325 4309 1202 ICV_9 $T=734080 487320 0 0 $X=734080 $Y=486940
X3624 4492 4415 2 1 4425 4459 4288 4281 4461 4480 3985 1202 ICV_9 $T=767560 447000 1 0 $X=767560 $Y=441580
X3625 4537 4356 2 1 4542 4550 4443 4433 4520 4527 4490 1202 ICV_9 $T=775620 376440 0 0 $X=775620 $Y=376060
X3626 4541 4426 2 1 4557 4459 4242 4271 4528 4533 3919 1202 ICV_9 $T=776860 467160 0 0 $X=776860 $Y=466780
X3627 4575 654 2 1 4587 662 653 655 4562 4548 4567 1202 ICV_9 $T=786160 527640 0 0 $X=786160 $Y=527260
X3628 4598 4385 2 1 4624 4610 4578 4530 4577 4535 4556 1202 ICV_9 $T=791740 436920 1 0 $X=791740 $Y=431500
X3629 4654 4430 2 1 4675 4597 4410 4412 4622 4646 675 1202 ICV_9 $T=802280 406680 1 0 $X=802280 $Y=401260
X3630 4655 4524 2 1 4669 4464 4635 4614 4603 4643 4612 1202 ICV_9 $T=802280 507480 1 0 $X=802280 $Y=502060
X3631 4697 4524 2 1 4709 4436 4635 4614 4657 4645 4690 1202 ICV_9 $T=809720 487320 0 0 $X=809720 $Y=486940
X3632 4701 4524 2 1 4713 4423 4635 4614 4679 3844 4698 1202 ICV_9 $T=811580 497400 0 0 $X=811580 $Y=497020
X3633 4702 629 2 1 4714 670 4667 655 4685 4694 4681 1202 ICV_9 $T=811580 527640 0 0 $X=811580 $Y=527260
X3634 4897 4898 2 1 4924 756 735 736 4880 4873 4892 1202 ICV_9 $T=855600 497400 0 0 $X=855600 $Y=497020
X3635 4879 763 2 1 768 722 750 744 4852 740 743 1202 ICV_9 $T=856220 537720 1 0 $X=856220 $Y=532300
X3636 4921 4898 2 1 4848 4917 4894 4903 4887 4905 4909 1202 ICV_9 $T=858700 467160 1 0 $X=858700 $Y=461740
X3637 4966 4951 2 1 5059 797 4875 4891 5016 802 4946 1202 ICV_9 $T=881020 376440 1 0 $X=881020 $Y=371020
X3638 5144 5092 2 1 5187 4695 5008 5084 5152 5110 5119 1202 ICV_9 $T=907680 477240 1 0 $X=907680 $Y=471820
X3639 5607 5603 2 1 5629 5554 5573 5477 5508 5587 5591 1202 ICV_9 $T=1001920 406680 1 0 $X=1001920 $Y=401260
X3640 5659 5466 2 1 5672 1023 5512 5519 5589 5648 5647 1202 ICV_9 $T=1013080 447000 0 0 $X=1013080 $Y=446620
X3641 5716 1020 2 1 5718 5554 1003 1030 5700 5692 5707 1202 ICV_9 $T=1026720 376440 0 0 $X=1026720 $Y=376060
X3642 1046 1042 2 1 1050 5554 991 5728 5708 5731 1045 1202 ICV_9 $T=1032300 366360 0 0 $X=1032300 $Y=365980
X3643 5757 980 2 1 5779 5668 1047 5728 5732 5739 5719 1202 ICV_9 $T=1036020 406680 1 0 $X=1036020 $Y=401260
X3644 5898 5854 2 1 5912 5895 5760 5680 5875 5782 5889 1202 ICV_9 $T=1065160 426840 1 0 $X=1065160 $Y=421420
X3645 1111 1084 2 1 5965 6027 1028 1087 5989 6013 1108 1202 ICV_9 $T=1093060 386520 1 0 $X=1093060 $Y=381100
X3646 6034 5881 2 1 6051 5907 6005 5816 5942 6020 1110 1202 ICV_9 $T=1094300 477240 1 0 $X=1094300 $Y=471820
X3647 6072 5881 2 1 6091 1123 6005 5816 6052 6045 1117 1202 ICV_9 $T=1102980 477240 1 0 $X=1102980 $Y=471820
X3648 5798 5836 2 1 6098 6099 1102 5966 6058 6063 5774 1202 ICV_9 $T=1103600 517560 0 0 $X=1103600 $Y=517180
X3649 6075 1083 2 1 6103 6043 1028 1087 5967 6054 6036 1202 ICV_9 $T=1104220 386520 1 0 $X=1104220 $Y=381100
X3650 6093 5842 2 1 6115 6099 6068 5829 6073 6085 6084 1202 ICV_9 $T=1106700 497400 1 0 $X=1106700 $Y=491980
X3651 6100 5880 2 1 6129 6074 6042 5973 6070 6087 6088 1202 ICV_9 $T=1107940 457080 1 0 $X=1107940 $Y=451660
X3652 2516 1 2 2549 2508 231 256 2380 1202 ICV_11 $T=442680 507480 0 0 $X=442680 $Y=507100
X3653 3919 1 2 3951 3957 3926 3986 3988 1202 ICV_11 $T=656580 477240 1 0 $X=656580 $Y=471820
X3654 3985 1 2 4001 4005 3926 4056 3990 1202 ICV_11 $T=667740 447000 1 0 $X=667740 $Y=441580
X3655 4013 1 2 4050 4049 3926 3981 3825 1202 ICV_11 $T=674560 477240 0 0 $X=674560 $Y=476860
X3656 4020 1 2 4047 4055 541 4056 4095 1202 ICV_11 $T=675180 416760 0 0 $X=675180 $Y=416380
X3657 4150 1 2 4126 4174 3926 4156 3804 1202 ICV_11 $T=698740 447000 0 0 $X=698740 $Y=446620
X3658 4229 1 2 4258 4259 3926 4303 4229 1202 ICV_11 $T=718580 436920 0 0 $X=718580 $Y=436540
X3659 4243 1 2 4269 4246 3926 4237 4243 1202 ICV_11 $T=720440 457080 1 0 $X=720440 $Y=451660
X3660 4419 1 2 4437 4442 612 4483 4505 1202 ICV_11 $T=756400 507480 0 0 $X=756400 $Y=507100
X3661 4535 1 2 4551 4545 628 4570 4506 1202 ICV_11 $T=778720 426840 1 0 $X=778720 $Y=421420
X3662 4952 1 2 4969 4979 4560 4935 5035 1202 ICV_11 $T=868620 487320 0 0 $X=868620 $Y=486940
X3663 837 1 2 842 5224 820 849 5257 1202 ICV_11 $T=916980 537720 1 0 $X=916980 $Y=532300
X3664 5227 1 2 5248 5252 820 5285 5227 1202 ICV_11 $T=922560 517560 1 0 $X=922560 $Y=512140
X3665 5624 1 2 5655 5673 943 5674 1033 1202 ICV_11 $T=1015560 517560 0 0 $X=1015560 $Y=517180
X3666 5692 1 2 5691 5718 1039 5751 5707 1202 ICV_11 $T=1025480 386520 1 0 $X=1025480 $Y=381100
X3667 5772 1 2 5776 5796 1039 5748 1075 1202 ICV_11 $T=1042840 457080 0 0 $X=1042840 $Y=456700
X3668 1081 1 2 1085 5878 1066 1091 5846 1202 ICV_11 $T=1060200 537720 1 0 $X=1060200 $Y=532300
X3669 5889 1 2 5898 5894 1039 5950 5782 1202 ICV_11 $T=1068880 426840 0 0 $X=1068880 $Y=426460
X3670 5920 1 2 5935 5953 1039 5990 5997 1202 ICV_11 $T=1076320 416760 1 0 $X=1076320 $Y=411340
X3671 3992 4022 2 1 3964 517 536 4002 4038 4015 3980 1202 ICV_13 $T=675800 457080 0 180 $X=671460 $Y=451660
X3672 4292 3995 2 1 4267 4228 4316 4306 4272 4300 4296 1202 ICV_13 $T=730360 507480 0 180 $X=726020 $Y=502060
X3673 4424 4382 2 1 4379 4399 4441 4216 4449 4420 3874 1202 ICV_13 $T=757640 497400 0 180 $X=753300 $Y=491980
X3674 640 615 2 1 639 637 642 575 4467 641 623 1202 ICV_13 $T=766320 366360 1 180 $X=761980 $Y=365980
X3675 4596 4430 2 1 4563 4518 4410 4412 4599 668 667 1202 ICV_13 $T=796080 406680 0 180 $X=791740 $Y=401260
X3676 4773 4776 2 1 4734 4737 4797 4790 4795 4733 4780 1202 ICV_13 $T=835140 477240 0 180 $X=830800 $Y=471820
X3677 4819 4822 2 1 4804 731 4872 4858 4866 4801 4744 1202 ICV_13 $T=850640 477240 0 180 $X=846300 $Y=471820
X3678 5058 4781 2 1 4979 5037 5008 4823 5070 5042 5035 1202 ICV_13 $T=890320 487320 1 180 $X=885980 $Y=486940
X3679 5072 4883 2 1 5044 797 5091 4933 5015 5071 5066 1202 ICV_13 $T=892800 406680 0 180 $X=888460 $Y=401260
X3680 5194 4841 2 1 5182 821 5089 4983 5231 5190 5174 1202 ICV_13 $T=921320 507480 1 180 $X=916980 $Y=507100
X3681 5559 980 2 1 5542 904 991 978 5580 5553 5537 1202 ICV_13 $T=998200 376440 0 180 $X=993860 $Y=371020
X3682 5696 5681 2 1 5678 1023 5709 5519 5712 5686 5650 1202 ICV_13 $T=1026100 447000 1 180 $X=1021760 $Y=446620
X3683 5873 1084 2 1 5803 5856 1028 1087 5892 5869 5850 1202 ICV_13 $T=1065160 386520 0 180 $X=1060820 $Y=381100
X3684 1086 1042 2 1 5802 5856 1059 1082 5886 1088 1078 1202 ICV_13 $T=1066400 366360 1 180 $X=1062060 $Y=365980
X3685 5862 5790 2 1 5808 5856 5754 5896 5871 5841 5860 1202 ICV_13 $T=1067020 396600 0 180 $X=1062680 $Y=391180
X3686 5916 5842 2 1 5903 5410 5749 5829 5933 5917 5901 1202 ICV_13 $T=1074460 497400 0 180 $X=1070120 $Y=491980
X3687 6035 5836 2 1 6017 5999 1102 5966 6049 5979 6041 1202 ICV_13 $T=1099260 517560 1 180 $X=1094920 $Y=517180
X3688 2581 1 2 2557 2517 231 2488 2581 1202 ICV_15 $T=442060 477240 0 0 $X=442060 $Y=476860
X3689 529 1 2 3991 3936 518 3972 3956 1202 ICV_15 $T=658440 527640 1 0 $X=658440 $Y=522220
X3690 4391 1 2 4370 4340 3926 4303 4391 1202 ICV_15 $T=739040 447000 0 0 $X=739040 $Y=446620
X3691 4656 1 2 4671 4608 4560 4539 4644 1202 ICV_15 $T=796700 457080 1 0 $X=796700 $Y=451660
X3692 4766 1 2 4765 4726 4560 4751 707 1202 ICV_15 $T=822120 447000 0 0 $X=822120 $Y=446620
X3693 4784 1 2 4771 4731 628 4756 713 1202 ICV_15 $T=824600 396600 1 0 $X=824600 $Y=391180
X3694 4780 1 2 4773 4734 4560 4768 4780 1202 ICV_15 $T=825840 487320 1 0 $X=825840 $Y=481900
X3695 4735 1 2 4736 4747 628 4756 4730 1202 ICV_15 $T=828940 376440 1 0 $X=828940 $Y=371020
X3696 4881 1 2 4906 4824 718 4756 4834 1202 ICV_15 $T=844440 386520 1 0 $X=844440 $Y=381100
X3697 4986 1 2 4963 4945 718 4893 4986 1202 ICV_15 $T=867380 416760 1 0 $X=867380 $Y=411340
X3698 5199 1 2 5205 5214 820 5236 5186 1202 ICV_15 $T=920080 426840 0 0 $X=920080 $Y=426460
X3699 5173 1 2 5162 5225 820 5261 863 1202 ICV_15 $T=923180 467160 0 0 $X=923180 $Y=466780
X3700 5211 1 2 5243 5245 718 5236 868 1202 ICV_15 $T=926900 396600 0 0 $X=926900 $Y=396220
X3701 5295 1 2 5324 5281 820 5285 5270 1202 ICV_15 $T=934340 497400 0 0 $X=934340 $Y=497020
X3702 5305 1 2 5315 5282 820 849 5305 1202 ICV_15 $T=934340 527640 0 0 $X=934340 $Y=527260
X3703 5587 1 2 5607 5550 846 5594 968 1202 ICV_15 $T=996340 396600 1 0 $X=996340 $Y=391180
X3704 5648 1 2 5616 5597 943 5348 5648 1202 ICV_15 $T=1004400 447000 1 0 $X=1004400 $Y=441580
X3705 5818 1 2 5855 5837 1039 5834 5870 1202 ICV_15 $T=1055860 416760 1 0 $X=1055860 $Y=411340
X3706 5948 1 2 5952 5923 1039 5957 5948 1202 ICV_15 $T=1075700 376440 0 0 $X=1075700 $Y=376060
X3707 6041 1 2 6035 5996 1066 1100 5983 1202 ICV_15 $T=1089960 527640 0 0 $X=1089960 $Y=527260
X3708 49 2 1386 1 1359 1396 1202 ICV_16 $T=253580 507480 1 0 $X=253580 $Y=502060
X3709 1656 2 1669 1 1668 1688 1202 ICV_16 $T=305660 396600 1 0 $X=305660 $Y=391180
X3710 1828 2 1894 1 1791 1902 1202 ICV_16 $T=341620 386520 1 0 $X=341620 $Y=381100
X3711 305 2 2547 1 305 2742 1202 ICV_16 $T=485460 477240 0 0 $X=485460 $Y=476860
X3712 2918 2 3014 1 2938 3026 1202 ICV_16 $T=517700 396600 0 0 $X=517700 $Y=396220
X3713 3067 2 3151 1 3139 378 1202 ICV_16 $T=533200 376440 0 0 $X=533200 $Y=376060
X3714 275 2 3226 1 3226 3115 1202 ICV_16 $T=543740 416760 0 0 $X=543740 $Y=416380
X3715 3548 2 3576 1 3463 3592 1202 ICV_16 $T=602020 396600 1 0 $X=602020 $Y=391180
X3716 3709 2 473 1 473 3760 1202 ICV_16 $T=626820 386520 0 0 $X=626820 $Y=386140
X3717 2465 2 4404 1 4418 4431 1202 ICV_16 $T=757640 447000 1 0 $X=757640 $Y=441580
X3718 4433 2 4398 1 4323 4446 1202 ICV_16 $T=760740 396600 0 0 $X=760740 $Y=396220
X3719 4398 2 4450 1 4446 4465 1202 ICV_16 $T=763220 396600 0 0 $X=763220 $Y=396220
X3720 4670 2 689 1 689 692 1202 ICV_16 $T=817160 366360 0 0 $X=817160 $Y=365980
X3721 4941 2 5146 1 5146 5153 1202 ICV_16 $T=906440 376440 0 0 $X=906440 $Y=376060
X3722 4695 2 5201 1 5201 5207 1202 ICV_16 $T=920080 477240 1 0 $X=920080 $Y=471820
X3723 5449 2 5457 1 5461 5466 1202 ICV_16 $T=977120 457080 0 0 $X=977120 $Y=456700
X3724 5489 2 5611 1 5611 5604 1202 ICV_16 $T=1005640 487320 0 0 $X=1005640 $Y=486940
X3725 208 1923 1 2 INV6CK $T=412300 477240 0 0 $X=412300 $Y=476860
X3726 951 954 1 2 INV6CK $T=982080 386520 0 0 $X=982080 $Y=386140
X3727 4593 4511 4632 4648 4661 1 2 AN4 $T=802280 396600 1 0 $X=802280 $Y=391180
X3728 5871 5875 5886 5892 5090 1 2 AN4 $T=1065780 386520 0 0 $X=1065780 $Y=386140
X3729 5943 5976 5940 5967 4982 1 2 AN4 $T=1088100 396600 0 180 $X=1081900 $Y=391180
X3730 6025 6049 6050 6039 5021 1 2 AN4 $T=1104220 497400 0 180 $X=1098020 $Y=491980
X3731 6073 6077 6070 6066 5185 1 2 AN4 $T=1109180 487320 1 180 $X=1102980 $Y=486940
X3732 19 1246 10 1 2 ND2 $T=230020 517560 1 0 $X=230020 $Y=512140
X3733 366 3179 378 1 2 ND2 $T=538780 386520 0 180 $X=536920 $Y=381100
X3734 3190 3207 3180 1 2 ND2 $T=540640 416760 1 0 $X=540640 $Y=411340
X3735 3215 3078 3207 1 2 ND2 $T=543120 406680 1 180 $X=541260 $Y=406300
X3736 3237 3239 3238 1 2 ND2 $T=546220 396600 1 0 $X=546220 $Y=391180
X3737 3249 3248 3213 1 2 ND2 $T=548080 376440 1 0 $X=548080 $Y=371020
X3738 3304 3299 2842 1 2 ND2 $T=556760 396600 1 180 $X=554900 $Y=396220
X3739 3320 3306 3296 1 2 ND2 $T=558620 386520 1 0 $X=558620 $Y=381100
X3740 3359 404 3361 1 2 ND2 $T=565440 376440 1 0 $X=565440 $Y=371020
X3741 3375 3334 3366 1 2 ND2 $T=569160 396600 0 180 $X=567300 $Y=391180
X3742 3387 3388 3360 1 2 ND2 $T=571020 396600 1 0 $X=571020 $Y=391180
X3743 3392 3393 3131 1 2 ND2 $T=572260 406680 1 0 $X=572260 $Y=401260
X3744 3399 3318 3412 1 2 ND2 $T=574120 406680 1 0 $X=574120 $Y=401260
X3745 3417 3222 3430 1 2 ND2 $T=575980 406680 0 0 $X=575980 $Y=406300
X3746 3414 3449 3382 1 2 ND2 $T=577840 436920 1 0 $X=577840 $Y=431500
X3747 3495 3445 3509 1 2 ND2 $T=588380 386520 0 0 $X=588380 $Y=386140
X3748 3521 3519 3528 1 2 ND2 $T=592100 406680 1 0 $X=592100 $Y=401260
X3749 3513 3533 3538 1 2 ND2 $T=593960 447000 0 0 $X=593960 $Y=446620
X3750 3541 3505 3532 1 2 ND2 $T=595820 426840 1 0 $X=595820 $Y=421420
X3751 3535 3545 3550 1 2 ND2 $T=595820 507480 0 0 $X=595820 $Y=507100
X3752 3533 3554 3506 1 2 ND2 $T=599540 447000 0 180 $X=597680 $Y=441580
X3753 3522 3549 3567 1 2 ND2 $T=598300 416760 0 0 $X=598300 $Y=416380
X3754 3690 3669 3672 1 2 ND2 $T=616900 436920 1 180 $X=615040 $Y=436540
X3755 3601 3715 3545 1 2 ND2 $T=620620 507480 1 180 $X=618760 $Y=507100
X3756 3723 3686 3692 1 2 ND2 $T=623720 426840 1 180 $X=621860 $Y=426460
X3757 3731 3537 3745 1 2 ND2 $T=623720 426840 0 0 $X=623720 $Y=426460
X3758 3772 3606 3793 1 2 ND2 $T=633020 436920 1 0 $X=633020 $Y=431500
X3759 3780 3773 3762 1 2 ND2 $T=633020 457080 1 0 $X=633020 $Y=451660
X3760 3800 3780 3791 1 2 ND2 $T=636740 447000 1 180 $X=634880 $Y=446620
X3761 3789 3791 3790 1 2 ND2 $T=636740 457080 0 180 $X=634880 $Y=451660
X3762 486 3818 479 1 2 ND2 $T=639840 537720 0 180 $X=637980 $Y=532300
X3763 3795 3819 3818 1 2 ND2 $T=641700 537720 0 180 $X=639840 $Y=532300
X3764 3819 3834 3832 1 2 ND2 $T=643560 517560 1 180 $X=641700 $Y=517180
X3765 3830 3843 3854 1 2 ND2 $T=644180 507480 0 0 $X=644180 $Y=507100
X3766 3867 3880 3888 1 2 ND2 $T=649760 487320 1 0 $X=649760 $Y=481900
X3767 3880 3879 3887 1 2 ND2 $T=650380 447000 0 0 $X=650380 $Y=446620
X3768 3843 3910 3866 1 2 ND2 $T=654720 467160 1 180 $X=652860 $Y=466780
X3769 506 3911 3900 1 2 ND2 $T=655960 507480 1 180 $X=654100 $Y=507100
X3770 3022 3050 2992 3067 2 1 2985 OA112 $T=521420 386520 1 0 $X=521420 $Y=381100
X3771 3121 3149 3106 3067 2 1 3152 OA112 $T=532580 416760 1 0 $X=532580 $Y=411340
X3772 3293 3300 3119 3310 2 1 3330 OA112 $T=554900 487320 0 0 $X=554900 $Y=486940
X3773 1923 114 1 2 INV8CK $T=347820 416760 0 180 $X=341000 $Y=411340
X3774 130 1886 1 133 1914 134 2 OAI112HS $T=342860 366360 0 0 $X=342860 $Y=365980
X3775 129 1915 1 1931 1936 1941 2 OAI112HS $T=345960 376440 1 0 $X=345960 $Y=371020
X3776 2684 2586 1 2714 2720 2723 2 OAI112HS $T=473060 487320 1 0 $X=473060 $Y=481900
X3777 2879 2992 1 2977 2944 2959 2 OAI112HS $T=517700 376440 1 180 $X=513360 $Y=376060
X3778 352 2954 1 2973 2910 2987 2 OAI112HS $T=518940 416760 1 180 $X=514600 $Y=416380
X3779 2879 3106 1 3060 3083 3079 2 OAI112HS $T=530720 416760 0 180 $X=526380 $Y=411340
X3780 2879 3133 1 3120 3110 3097 2 OAI112HS $T=533200 386520 1 180 $X=528860 $Y=386140
X3781 3067 3133 1 3179 3201 3170 2 OAI112HS $T=536920 386520 0 0 $X=536920 $Y=386140
X3782 1209 10 2 19 1238 1209 1 AOI22H $T=220720 517560 1 0 $X=220720 $Y=512140
X3783 4621 792 4982 4985 1 2 ND3P $T=872340 396600 1 0 $X=872340 $Y=391180
X3784 4649 789 5005 4901 1 2 ND3P $T=881020 396600 1 180 $X=876060 $Y=396220
X3785 4477 799 5009 5012 1 2 ND3P $T=877300 406680 1 0 $X=877300 $Y=401260
X3786 4674 828 5165 5161 1 2 ND3P $T=914500 487320 1 180 $X=909540 $Y=486940
X3787 3376 2 3389 1 3243 NR2P $T=571640 416760 0 180 $X=567920 $Y=411340
X3788 1902 1894 1915 2 129 1 1922 AN4B1S $T=344100 386520 1 0 $X=344100 $Y=381100
X3789 1959 151 2011 2 153 1 2000 AN4B1S $T=357740 376440 1 0 $X=357740 $Y=371020
X3790 2000 1921 1918 2 2016 1 2025 AN4B1S $T=357740 386520 1 0 $X=357740 $Y=381100
X3791 2401 2405 213 2 216 1 2400 AN4B1S $T=425940 376440 0 180 $X=421600 $Y=371020
X3792 2420 223 2095 2 1845 1 2401 AN4B1S $T=427800 386520 0 180 $X=423460 $Y=381100
X3793 3101 368 3086 2 3058 1 3087 AN4B1S $T=528860 376440 0 180 $X=524520 $Y=371020
X3794 3277 3144 3264 2 3258 1 3241 AN4B1S $T=553040 386520 1 180 $X=548700 $Y=386140
X3795 4148 4140 4141 2 4081 1 559 AN4B1S $T=700600 497400 1 180 $X=696260 $Y=497020
X3796 4122 4124 4142 2 4149 1 560 AN4B1S $T=696260 537720 1 0 $X=696260 $Y=532300
X3797 4155 4112 4167 2 4100 1 567 AN4B1S $T=700600 497400 0 0 $X=700600 $Y=497020
X3798 4208 4203 4200 2 4194 1 573 AN4B1S $T=713000 497400 1 180 $X=708660 $Y=497020
X3799 4211 4170 4202 2 4115 1 577 AN4B1S $T=713620 426840 0 180 $X=709280 $Y=421420
X3800 4199 4182 4204 2 4121 1 580 AN4B1S $T=709900 416760 0 0 $X=709900 $Y=416380
X3801 4313 4310 4305 2 4298 1 590 AN4B1S $T=734700 406680 1 180 $X=730360 $Y=406300
X3802 5463 5451 5358 2 5450 1 4202 AN4B1S $T=979600 396600 0 180 $X=975260 $Y=391180
X3803 5464 5452 5326 2 936 1 4305 AN4B1S $T=979600 396600 1 180 $X=975260 $Y=396220
X3804 5478 5484 5382 2 959 1 4204 AN4B1S $T=982080 406680 1 0 $X=982080 $Y=401260
X3805 5520 5498 5362 2 5506 1 4167 AN4B1S $T=990760 497400 1 180 $X=986420 $Y=497020
X3806 5548 5543 5353 2 5535 1 4200 AN4B1S $T=995720 487320 1 180 $X=991380 $Y=486940
X3807 5595 5582 5291 2 5578 1 4184 AN4B1S $T=1005020 416760 1 180 $X=1000680 $Y=416380
X3808 5625 5593 5367 2 5583 1 4142 AN4B1S $T=1006260 487320 0 180 $X=1001920 $Y=481900
X3809 5320 1 2 877 BUF3CK $T=942400 396600 1 0 $X=942400 $Y=391180
X3810 1300 2 1266 31 1306 1 1352 FA1S $T=233120 396600 1 0 $X=233120 $Y=391180
X3811 1315 2 1285 1248 1298 1 1354 FA1S $T=235600 396600 0 0 $X=235600 $Y=396220
X3812 36 2 1315 1344 1300 1 1356 FA1S $T=236220 386520 0 0 $X=236220 $Y=386140
X3813 1332 2 1329 34 1336 1 1344 FA1S $T=238080 376440 1 0 $X=238080 $Y=371020
X3814 1340 2 1335 1284 1312 1 1374 FA1S $T=239940 406680 1 0 $X=239940 $Y=401260
X3815 1376 2 1377 55 1332 1 42 FA1S $T=257300 366360 1 180 $X=245520 $Y=365980
X3816 1369 2 1303 1318 1388 1 1477 FA1S $T=246760 447000 1 0 $X=246760 $Y=441580
X3817 1377 2 1379 1358 1347 1 1411 FA1S $T=248620 416760 0 0 $X=248620 $Y=416380
X3818 1402 2 1373 1324 1430 1 1441 FA1S $T=253580 487320 1 0 $X=253580 $Y=481900
X3819 1406 2 1263 1423 1412 1 1443 FA1S $T=254200 426840 1 0 $X=254200 $Y=421420
X3820 1407 2 1398 1261 1380 1 1440 FA1S $T=254200 436920 0 0 $X=254200 $Y=436540
X3821 1416 2 1334 1273 1364 1 1454 FA1S $T=256060 426840 0 0 $X=256060 $Y=426460
X3822 1425 2 1357 1410 1418 1 1461 FA1S $T=258540 436920 1 0 $X=258540 $Y=431500
X3823 1426 2 1449 1270 1400 1 1468 FA1S $T=258540 457080 1 0 $X=258540 $Y=451660
X3824 1437 2 1411 1429 1356 1 1473 FA1S $T=261020 396600 1 0 $X=261020 $Y=391180
X3825 1438 2 1275 1424 1415 1 1474 FA1S $T=261020 447000 0 0 $X=261020 $Y=446620
X3826 1429 2 1425 1352 1340 1 1480 FA1S $T=262260 406680 1 0 $X=262260 $Y=401260
X3827 1460 2 1461 1483 1467 1 1422 FA1S $T=274660 416760 1 180 $X=262880 $Y=416380
X3828 1447 2 1271 1350 1455 1 1479 FA1S $T=262880 467160 1 0 $X=262880 $Y=461740
X3829 1452 2 1402 1468 1447 1 1489 FA1S $T=264120 457080 0 0 $X=264120 $Y=456700
X3830 1448 2 1416 1374 1406 1 1467 FA1S $T=264740 406680 0 0 $X=264740 $Y=406300
X3831 1459 2 1354 1448 1480 1 1504 FA1S $T=265360 396600 0 0 $X=265360 $Y=396220
X3832 69 2 1401 1339 1409 1 1503 FA1S $T=266600 376440 0 0 $X=266600 $Y=376060
X3833 1466 2 1369 1440 1438 1 1498 FA1S $T=267220 436920 0 0 $X=267220 $Y=436540
X3834 1476 2 1454 1466 1515 1 1520 FA1S $T=268460 426840 1 0 $X=268460 $Y=421420
X3835 1478 2 1342 1465 1475 1 1511 FA1S $T=269700 467160 0 0 $X=269700 $Y=466780
X3836 1483 2 1478 1443 1407 1 1515 FA1S $T=270320 426840 0 0 $X=270320 $Y=426460
X3837 1484 2 1518 1474 1426 1 1527 FA1S $T=271560 457080 1 0 $X=271560 $Y=451660
X3838 1490 2 1511 1484 1498 1 1529 FA1S $T=272800 436920 1 0 $X=272800 $Y=431500
X3839 72 2 1503 1376 74 1 78 FA1S $T=273420 366360 0 0 $X=273420 $Y=365980
X3840 1494 2 1451 1404 1487 1 1554 FA1S $T=273420 507480 1 0 $X=273420 $Y=502060
X3841 1502 2 1477 1452 1527 1 1536 FA1S $T=274660 447000 1 0 $X=274660 $Y=441580
X3842 1512 2 1494 1532 1513 1 1553 FA1S $T=275900 487320 1 0 $X=275900 $Y=481900
X3843 1496 2 1524 1304 1439 1 1532 FA1S $T=275900 487320 0 0 $X=275900 $Y=486940
X3844 1513 2 1292 1333 1506 1 1545 FA1S $T=275900 497400 1 0 $X=275900 $Y=491980
X3845 1517 2 1510 1501 1542 1 1548 FA1S $T=276520 406680 0 0 $X=276520 $Y=406300
X3846 1507 2 1528 1479 1496 1 1544 FA1S $T=276520 467160 1 0 $X=276520 $Y=461740
X3847 1521 2 1535 1507 1489 1 1540 FA1S $T=277760 457080 0 0 $X=277760 $Y=456700
X3848 1518 2 1381 1491 1508 1 1535 FA1S $T=278380 477240 1 0 $X=278380 $Y=471820
X3849 77 2 1495 1471 1555 1 1561 FA1S $T=279000 376440 1 0 $X=279000 $Y=371020
X3850 1541 2 1581 1562 1530 1 1509 FA1S $T=292020 386520 0 180 $X=280240 $Y=381100
X3851 1530 2 1497 1519 1565 1 1567 FA1S $T=280240 396600 1 0 $X=280240 $Y=391180
X3852 1546 2 1576 1561 1537 1 1516 FA1S $T=292640 376440 1 180 $X=280860 $Y=376060
X3853 1537 2 1514 1500 1571 1 1562 FA1S $T=281480 386520 0 0 $X=281480 $Y=386140
X3854 1528 2 1450 89 1538 1 1593 FA1S $T=283340 497400 0 0 $X=283340 $Y=497020
X3855 1549 2 1531 1533 1582 1 1589 FA1S $T=283960 416760 1 0 $X=283960 $Y=411340
X3856 1550 2 1441 1512 1544 1 1583 FA1S $T=283960 467160 0 0 $X=283960 $Y=466780
X3857 1556 2 1543 1539 1608 1 1603 FA1S $T=285200 426840 0 0 $X=285200 $Y=426460
X3858 1558 2 1587 1517 1567 1 1613 FA1S $T=285820 406680 1 0 $X=285820 $Y=401260
X3859 1559 2 1526 1586 1595 1 1601 FA1S $T=285820 416760 0 0 $X=285820 $Y=416380
X3860 1564 2 93 1362 1492 1 1617 FA1S $T=286440 507480 0 0 $X=286440 $Y=507100
X3861 1568 2 87 1463 1580 1 1618 FA1S $T=287060 527640 1 0 $X=287060 $Y=522220
X3862 1579 2 1551 1566 1557 1 1627 FA1S $T=288920 447000 0 0 $X=288920 $Y=446620
X3863 1566 2 1596 1552 1575 1 1624 FA1S $T=288920 457080 1 0 $X=288920 $Y=451660
X3864 1569 2 1577 1614 1609 1 1557 FA1S $T=301320 447000 0 180 $X=289540 $Y=441580
X3865 1563 2 1593 1570 1553 1 1628 FA1S $T=289540 487320 1 0 $X=289540 $Y=481900
X3866 1584 2 1619 1548 1549 1 1633 FA1S $T=290160 406680 0 0 $X=290160 $Y=406300
X3867 1599 2 1622 1569 1603 1 1560 FA1S $T=301940 426840 0 180 $X=290160 $Y=421420
X3868 1572 2 1554 1573 1630 1 1592 FA1S $T=290160 487320 0 0 $X=290160 $Y=486940
X3869 1570 2 94 1545 1564 1 1630 FA1S $T=290160 497400 1 0 $X=290160 $Y=491980
X3870 1573 2 1568 1617 1600 1 1643 FA1S $T=291400 507480 1 0 $X=291400 $Y=502060
X3871 1600 2 1393 1419 100 1 1647 FA1S $T=292640 517560 0 0 $X=292640 $Y=517180
X3872 1631 2 1672 1615 1624 1 1692 FA1S $T=296980 457080 0 0 $X=296980 $Y=456700
X3873 1615 2 1673 1588 1616 1 1693 FA1S $T=296980 467160 0 0 $X=296980 $Y=466780
X3874 1632 2 99 1427 1594 1 1714 FA1S $T=296980 527640 0 0 $X=296980 $Y=527260
X3875 1637 2 1681 1589 1559 1 1713 FA1S $T=297600 416760 1 0 $X=297600 $Y=411340
X3876 1648 2 1695 1685 1639 1 1605 FA1S $T=309380 497400 1 180 $X=297600 $Y=497020
X3877 1652 2 1698 1601 1556 1 1686 FA1S $T=299460 416760 0 0 $X=299460 $Y=416380
X3878 1653 2 102 1664 1643 1 1708 FA1S $T=299460 507480 0 0 $X=299460 $Y=507100
X3879 1682 2 103 104 101 1 1625 FA1S $T=311860 537720 0 180 $X=300080 $Y=532300
X3880 1664 2 1682 1647 1632 1 1724 FA1S $T=300700 527640 1 0 $X=300700 $Y=522220
X3881 1700 2 1736 1726 1604 1 1639 FA1S $T=313720 477240 1 180 $X=301940 $Y=476860
X3882 1707 2 1743 1700 1693 1 1642 FA1S $T=314340 477240 0 180 $X=302560 $Y=471820
X3883 1717 2 1618 1757 1724 1 1774 FA1S $T=306280 517560 0 0 $X=306280 $Y=517180
X3884 1750 2 1597 1470 1741 1 1800 FA1S $T=310620 527640 0 0 $X=310620 $Y=527260
X3885 1685 2 1802 1794 1725 1 1728 FA1S $T=324260 507480 0 180 $X=312480 $Y=502060
X3886 1757 2 113 1625 1714 1 1830 FA1S $T=314960 527640 1 0 $X=314960 $Y=522220
X3887 1747 2 1769 1814 1728 1 1825 FA1S $T=316200 507480 0 0 $X=316200 $Y=507100
X3888 1818 2 1849 1855 1829 1 1720 FA1S $T=331080 447000 0 180 $X=319300 $Y=441580
X3889 1819 2 120 115 1789 1 1856 FA1S $T=321780 537720 1 0 $X=321780 $Y=532300
X3890 1826 2 1819 121 1800 1 1863 FA1S $T=323020 527640 0 0 $X=323020 $Y=527260
X3891 1823 2 1834 1865 1861 1 1756 FA1S $T=337900 457080 1 180 $X=326120 $Y=456700
X3892 1852 2 1874 1999 1864 1 1824 FA1S $T=339140 477240 0 180 $X=327360 $Y=471820
X3893 1821 2 1750 1826 1830 1 1893 FA1S $T=328600 527640 1 0 $X=328600 $Y=522220
X3894 1814 2 1875 1940 1798 1 1838 FA1S $T=341000 507480 0 180 $X=329220 $Y=502060
X3895 1832 2 1833 1838 1883 1 1885 FA1S $T=329220 517560 1 0 $X=329220 $Y=512140
X3896 1858 2 119 1876 1863 1 1884 FA1S $T=329220 517560 0 0 $X=329220 $Y=517180
X3897 1870 2 1901 1851 1848 1 1834 FA1S $T=342240 457080 0 180 $X=330460 $Y=451660
X3898 1831 2 1889 1852 1873 1 1740 FA1S $T=342240 467160 0 180 $X=330460 $Y=461740
X3899 1857 2 1903 1879 1868 1 1748 FA1S $T=344100 436920 0 180 $X=332320 $Y=431500
X3900 1879 2 1904 1910 1870 1 1855 FA1S $T=344720 447000 0 180 $X=332940 $Y=441580
X3901 1829 2 1951 1905 1900 1 1861 FA1S $T=345960 447000 1 180 $X=334180 $Y=446620
X3902 1876 2 123 1856 127 1 1927 FA1S $T=335420 537720 1 0 $X=335420 $Y=532300
X3903 1899 2 1935 1909 1916 1 1868 FA1S $T=348440 426840 1 180 $X=336660 $Y=426460
X3904 1887 2 1574 1499 1926 1 1930 FA1S $T=336660 527640 0 0 $X=336660 $Y=527260
X3905 1877 2 1939 1899 1895 1 1723 FA1S $T=349060 426840 0 180 $X=337280 $Y=421420
X3906 1854 2 1934 1932 1824 1 1847 FA1S $T=350920 477240 1 180 $X=339140 $Y=476860
X3907 1901 2 1946 1958 1928 1 1880 FA1S $T=351540 457080 1 180 $X=339760 $Y=456700
X3908 1929 2 1957 1953 1938 1 1864 FA1S $T=352780 467160 1 180 $X=341000 $Y=466780
X3909 1937 2 1961 1984 1943 1 1895 FA1S $T=354020 416760 1 180 $X=342240 $Y=416380
X3910 1932 2 1963 1962 1947 1 1896 FA1S $T=354020 487320 0 180 $X=342240 $Y=481900
X3911 1938 2 1968 1964 1948 1 1897 FA1S $T=354020 487320 1 180 $X=342240 $Y=486940
X3912 1925 2 1887 132 1971 1 1978 FA1S $T=342860 527640 1 0 $X=342860 $Y=522220
X3913 1865 2 1880 1988 1929 1 1873 FA1S $T=355880 467160 0 180 $X=344100 $Y=461740
X3914 1841 2 1897 2004 1896 1 1881 FA1S $T=355880 497400 0 180 $X=344100 $Y=491980
X3915 1945 2 1981 1993 1966 1 1848 FA1S $T=356500 457080 0 180 $X=344720 $Y=451660
X3916 1961 2 1983 1977 1944 1 1909 FA1S $T=357120 436920 0 180 $X=345340 $Y=431500
X3917 1916 2 1945 1987 1950 1 1849 FA1S $T=358360 447000 0 180 $X=346580 $Y=441580
X3918 1883 2 2008 1994 1924 1 1919 FA1S $T=358360 517560 0 180 $X=346580 $Y=512140
X3919 1872 2 2012 1974 1985 1 1788 FA1S $T=358980 396600 0 180 $X=347200 $Y=391180
X3920 1907 2 2001 2013 1920 1 1775 FA1S $T=358980 406680 1 180 $X=347200 $Y=406300
X3921 1974 2 1954 2021 1986 1 1920 FA1S $T=359600 396600 1 180 $X=347820 $Y=396220
X3922 1878 2 2005 1937 1992 1 1733 FA1S $T=359600 416760 0 180 $X=347820 $Y=411340
X3923 1971 2 2010 1930 142 1 2031 FA1S $T=349680 527640 0 0 $X=349680 $Y=527260
X3924 1991 2 2017 2042 2002 1 1950 FA1S $T=362700 426840 1 180 $X=350920 $Y=426460
X3925 2002 2 2018 2030 2009 1 1951 FA1S $T=362700 447000 1 180 $X=350920 $Y=446620
X3926 1939 2 2041 2054 1991 1 1903 FA1S $T=363320 426840 0 180 $X=351540 $Y=421420
X3927 1999 2 2007 2022 2020 1 1962 FA1S $T=363940 477240 1 180 $X=352160 $Y=476860
X3928 1955 2 1997 2028 2006 1 1970 FA1S $T=365180 497400 1 180 $X=353400 $Y=497020
X3929 1898 2 1976 1919 2050 1 2056 FA1S $T=355260 517560 0 0 $X=355260 $Y=517180
X3930 2024 2 2065 2082 2035 1 1984 FA1S $T=367660 416760 1 180 $X=355880 $Y=416380
X3931 1839 2 2071 2039 2048 1 1780 FA1S $T=368900 376440 1 180 $X=357120 $Y=376060
X3932 1900 2 2059 2040 2055 1 1889 FA1S $T=369520 457080 1 180 $X=357740 $Y=456700
X3933 2040 2 2066 2060 2043 1 1874 FA1S $T=369520 467160 0 180 $X=357740 $Y=461740
X3934 1947 2 2069 2077 1996 1 1997 FA1S $T=370140 487320 0 180 $X=358360 $Y=481900
X3935 2004 2 2088 2087 2053 1 2006 FA1S $T=370140 497400 0 180 $X=358360 $Y=491980
X3936 2052 2 2084 2024 2064 1 1992 FA1S $T=371380 416760 0 180 $X=359600 $Y=411340
X3937 1977 2 2036 2094 2072 1 1904 FA1S $T=372000 436920 1 180 $X=360220 $Y=436540
X3938 2048 2 2103 2026 2075 1 1985 FA1S $T=372620 396600 0 180 $X=360840 $Y=391180
X3939 1908 2 2105 2052 2076 1 1732 FA1S $T=372620 406680 1 180 $X=360840 $Y=406300
X3940 2063 2 2113 2121 2081 1 2026 FA1S $T=373240 386520 1 180 $X=361460 $Y=386140
X3941 2068 2 2104 2114 2078 1 2021 FA1S $T=373860 406680 0 180 $X=362080 $Y=401260
X3942 1867 2 2115 164 2089 1 1770 FA1S $T=375720 366360 1 180 $X=363940 $Y=365980
X3943 2010 2 157 1525 2044 1 2120 FA1S $T=363940 527640 0 0 $X=363940 $Y=527260
X3944 2089 2 2063 2102 2090 1 2039 FA1S $T=376340 376440 0 180 $X=364560 $Y=371020
X3945 2065 2 2058 2129 2097 1 1935 FA1S $T=376340 426840 1 180 $X=364560 $Y=426460
X3946 2090 2 2118 2137 2068 1 2012 FA1S $T=376960 386520 0 180 $X=365180 $Y=381100
X3947 2082 2 2079 2140 2110 1 2054 FA1S $T=378200 426840 0 180 $X=366420 $Y=421420
X3948 1987 2 2135 2141 2125 1 1905 FA1S $T=379440 447000 0 180 $X=367660 $Y=441580
X3949 2050 2 2131 2083 1956 1 2147 FA1S $T=368280 517560 1 0 $X=368280 $Y=512140
X3950 1963 2 2142 2122 2133 1 2053 FA1S $T=380680 487320 1 180 $X=368900 $Y=486940
X3951 2107 2 2101 161 2120 1 2112 FA1S $T=369520 527640 1 0 $X=369520 $Y=522220
X3952 2101 2 160 159 163 1 2154 FA1S $T=369520 537720 1 0 $X=369520 $Y=532300
X3953 2084 2 2157 2172 2134 1 1943 FA1S $T=381920 416760 1 180 $X=370140 $Y=416380
X3954 1988 2 2150 2136 2138 1 1934 FA1S $T=381920 467160 0 180 $X=370140 $Y=461740
X3955 2047 2 2139 2027 2147 1 2165 FA1S $T=370760 507480 0 0 $X=370760 $Y=507100
X3956 2123 2 2176 2155 2143 1 2005 FA1S $T=383780 416760 0 180 $X=372000 $Y=411340
X3957 2087 2 2164 2159 2151 1 2099 FA1S $T=384400 497400 0 180 $X=372620 $Y=491980
X3958 2144 2 2099 2211 2116 1 2100 FA1S $T=385020 507480 0 180 $X=373240 $Y=502060
X3959 2013 2 2170 2123 2160 1 2076 FA1S $T=386260 406680 1 180 $X=374480 $Y=406300
X3960 2148 2 2132 2201 2173 1 2103 FA1S $T=386880 376440 1 180 $X=375100 $Y=376060
X3961 2121 2 2192 2191 2167 1 2114 FA1S $T=386880 396600 0 180 $X=375100 $Y=391180
X3962 2028 2 2183 2174 2169 1 2116 FA1S $T=386880 477240 0 180 $X=375100 $Y=471820
X3963 2166 2 2210 2175 2179 1 2081 FA1S $T=388120 386520 1 180 $X=376340 $Y=386140
X3964 2132 2 166 2215 2180 1 2104 FA1S $T=388120 396600 1 180 $X=376340 $Y=396220
X3965 170 2 175 2166 2185 1 2126 FA1S $T=388740 366360 1 180 $X=376960 $Y=365980
X3966 2115 2 165 2126 2148 1 2071 FA1S $T=377580 376440 1 0 $X=377580 $Y=371020
X3967 2161 2 2067 168 2154 1 2209 FA1S $T=378200 527640 0 0 $X=378200 $Y=527260
X3968 2113 2 2207 2204 2189 1 2078 FA1S $T=390600 386520 0 180 $X=378820 $Y=381100
X3969 1944 2 2162 2205 2177 1 1910 FA1S $T=391220 447000 0 180 $X=379440 $Y=441580
X3970 2171 2 2051 2203 2152 1 2229 FA1S $T=379440 517560 0 0 $X=379440 $Y=517180
X3971 1851 2 2156 2158 2163 1 2055 FA1S $T=380680 457080 0 0 $X=380680 $Y=456700
X3972 2139 2 2178 2197 2093 1 2152 FA1S $T=393080 517560 0 180 $X=381300 $Y=512140
X3973 2176 2 2230 2231 2223 1 2172 FA1S $T=395560 416760 1 180 $X=383780 $Y=416380
X3974 2035 2 2237 2232 2226 1 2041 FA1S $T=395560 426840 0 180 $X=383780 $Y=421420
X3975 2200 2 169 172 177 1 2249 FA1S $T=383780 537720 1 0 $X=383780 $Y=532300
X3976 2169 2 2263 2206 2228 1 2195 FA1S $T=399280 467160 1 180 $X=387500 $Y=466780
X3977 2211 2 2208 2109 2196 1 2258 FA1S $T=387500 487320 1 0 $X=387500 $Y=481900
X3978 2243 2 2266 2258 2195 1 2199 FA1S $T=399900 477240 0 180 $X=388120 $Y=471820
X3979 189 2 2250 2285 191 1 2102 FA1S $T=401760 366360 1 180 $X=389980 $Y=365980
X3980 2185 2 2273 2286 2262 1 2118 FA1S $T=401760 376440 0 180 $X=389980 $Y=371020
X3981 2250 2 2252 2281 2241 1 2173 FA1S $T=401760 376440 1 180 $X=389980 $Y=376060
X3982 2203 2 2295 2278 2214 1 2218 FA1S $T=402380 527640 0 180 $X=390600 $Y=522220
X3983 2257 2 2074 2240 2218 1 2314 FA1S $T=393700 517560 0 0 $X=393700 $Y=517180
X3984 2265 2 2244 2234 2259 1 2305 FA1S $T=394940 396600 1 0 $X=394940 $Y=391180
X3985 1986 2 2305 2313 2303 1 2160 FA1S $T=409200 406680 0 180 $X=397420 $Y=401260
X3986 2289 2 2254 2247 2315 1 2322 FA1S $T=398040 406680 0 0 $X=398040 $Y=406300
X3987 2170 2 2322 2316 2307 1 2064 FA1S $T=410440 416760 0 180 $X=398660 $Y=411340
X3988 2302 2 2312 2326 2274 1 2313 FA1S $T=401140 386520 0 0 $X=401140 $Y=386140
X3989 2307 2 2272 2327 2337 1 2134 FA1S $T=413540 416760 1 180 $X=401760 $Y=416380
X3990 2308 2 2296 2276 2287 1 2157 FA1S $T=402380 436920 1 0 $X=402380 $Y=431500
X3991 2323 2 2351 2338 2342 1 2284 FA1S $T=414160 497400 0 180 $X=402380 $Y=491980
X3992 2311 2 2332 2294 2297 1 2354 FA1S $T=402380 507480 0 0 $X=402380 $Y=507100
X3993 2319 2 2124 2304 2311 1 2359 FA1S $T=403620 517560 1 0 $X=403620 $Y=512140
X3994 2266 2 2310 2291 2329 1 2371 FA1S $T=407340 467160 1 0 $X=407340 $Y=461740
X3995 2240 2 2346 2387 2261 1 2304 FA1S $T=420360 517560 1 180 $X=408580 $Y=517180
X3996 2353 2 2330 2331 2382 1 2385 FA1S $T=409200 467160 0 0 $X=409200 $Y=466780
X3997 209 2 199 2340 2325 1 2285 FA1S $T=409820 376440 1 0 $X=409820 $Y=371020
X3998 2356 2 2301 2324 2308 1 2143 FA1S $T=409820 447000 0 0 $X=409820 $Y=446620
X3999 2201 2 2321 2300 2355 1 2392 FA1S $T=411060 376440 0 0 $X=411060 $Y=376060
X4000 2364 2 2368 2343 211 1 219 FA1S $T=411060 537720 1 0 $X=411060 $Y=532300
X4001 2369 2 2335 2348 2362 1 2388 FA1S $T=412300 416760 1 0 $X=412300 $Y=411340
X4002 2137 2 2265 2302 2392 1 2397 FA1S $T=412920 386520 0 0 $X=412920 $Y=386140
X4003 2075 2 2369 2393 2397 1 2001 FA1S $T=425320 396600 0 180 $X=413540 $Y=391180
X4004 2373 2 2345 2328 2357 1 2382 FA1S $T=413540 457080 1 0 $X=413540 $Y=451660
X4005 1954 2 2378 2381 2356 1 2105 FA1S $T=414780 426840 0 0 $X=414780 $Y=426460
X4006 2379 2 2309 2371 2373 1 2283 FA1S $T=414780 457080 0 0 $X=414780 $Y=456700
X4007 2393 2 2398 2289 2388 1 2303 FA1S $T=427180 406680 0 180 $X=415400 $Y=401260
X4008 2378 2 2306 2350 2367 1 2316 FA1S $T=415400 426840 1 0 $X=415400 $Y=421420
X4009 2381 2 2275 2336 2370 1 2155 FA1S $T=415400 436920 1 0 $X=415400 $Y=431500
X4010 2389 2 2365 2366 2406 1 2384 FA1S $T=417880 487320 0 0 $X=417880 $Y=486940
X4011 2395 2 2396 2333 2354 1 2459 FA1S $T=417880 517560 1 0 $X=417880 $Y=512140
X4012 2396 2 2360 2376 2279 1 2434 FA1S $T=417880 527640 1 0 $X=417880 $Y=522220
X4013 2404 2 2358 2391 214 1 2445 FA1S $T=419740 527640 0 0 $X=419740 $Y=527260
X4014 2431 2 2404 2339 2434 1 2458 FA1S $T=424080 517560 0 0 $X=424080 $Y=517180
X4015 2435 2 2364 221 2445 1 2474 FA1S $T=424700 537720 1 0 $X=424700 $Y=532300
X4016 2482 2 2515 2503 2460 1 2452 FA1S $T=444540 436920 1 180 $X=432760 $Y=436540
X4017 2481 2 2512 2447 2513 1 2532 FA1S $T=433380 386520 1 0 $X=433380 $Y=381100
X4018 2493 2 2466 2425 2486 1 2545 FA1S $T=435240 406680 0 0 $X=435240 $Y=406300
X4019 251 2 2471 2502 2481 1 2566 FA1S $T=439580 376440 1 0 $X=439580 $Y=371020
X4020 2541 2 2498 2509 2550 1 2487 FA1S $T=451360 416760 1 180 $X=439580 $Y=416380
X4021 2534 2 2522 2524 2493 1 2577 FA1S $T=441440 396600 0 0 $X=441440 $Y=396220
X4022 2588 2 2548 2545 2598 1 2609 FA1S $T=450740 406680 0 0 $X=450740 $Y=406300
X4023 2591 2 2559 2532 2602 1 2636 FA1S $T=451360 376440 0 0 $X=451360 $Y=376060
X4024 6142 2 2644 2651 2635 1 2580 FA1S $T=465000 517560 1 180 $X=453220 $Y=517180
X4025 2612 2 2597 2566 2591 1 2660 FA1S $T=455080 376440 1 0 $X=455080 $Y=371020
X4026 2642 2 2639 2614 2577 1 2643 FA1S $T=459420 396600 0 0 $X=459420 $Y=396220
X4027 2697 2 293 2681 2660 1 2711 FA1S $T=468720 376440 1 0 $X=468720 $Y=371020
X4028 294 2 292 2612 291 1 2772 FA1S $T=474300 366360 0 0 $X=474300 $Y=365980
X4029 2716 2 2534 2713 2636 1 2702 FA1S $T=474920 386520 0 0 $X=474920 $Y=386140
X4030 6143 2 335 325 330 1 2819 FA1S $T=509020 537720 0 180 $X=497240 $Y=532300
X4031 2881 2 2846 2863 2903 1 2951 FA1S $T=498480 477240 1 0 $X=498480 $Y=471820
X4032 2889 2 2859 2862 2881 1 2946 FA1S $T=499100 487320 1 0 $X=499100 $Y=481900
X4033 2903 2 2878 2887 2950 1 2980 FA1S $T=502200 467160 0 0 $X=502200 $Y=466780
X4034 2925 2 2877 2897 2889 1 2990 FA1S $T=504060 487320 0 0 $X=504060 $Y=486940
X4035 2931 2 2924 2964 2979 1 2999 FA1S $T=504680 457080 1 0 $X=504680 $Y=451660
X4036 2950 2 2865 2961 2931 1 3044 FA1S $T=510260 467160 1 0 $X=510260 $Y=461740
X4037 3004 2 3039 2955 3040 1 3055 FA1S $T=512120 477240 1 0 $X=512120 $Y=471820
X4038 3005 2 2898 2981 2925 1 3070 FA1S $T=512120 487320 1 0 $X=512120 $Y=481900
X4039 3017 2 2975 3027 3028 1 3069 FA1S $T=513360 457080 0 0 $X=513360 $Y=456700
X4040 3028 2 2896 3003 3004 1 3091 FA1S $T=515220 467160 0 0 $X=515220 $Y=466780
X4041 3040 2 3065 3016 3005 1 3105 FA1S $T=517080 477240 0 0 $X=517080 $Y=476860
X4042 3099 2 2876 3063 3088 1 3161 FA1S $T=523280 436920 0 0 $X=523280 $Y=436540
X4043 3116 2 2902 3075 3099 1 3112 FA1S $T=525140 447000 0 0 $X=525140 $Y=446620
X4044 2979 2 2893 3130 3116 1 3208 FA1S $T=528240 457080 1 0 $X=528240 $Y=451660
X4045 3255 2 3290 3308 3259 1 3216 FA1S $T=554280 457080 1 180 $X=542500 $Y=456700
X4046 3343 2 3357 3302 3353 1 3294 FA1S $T=567920 457080 1 180 $X=556140 $Y=456700
X4047 3328 2 3400 3343 3380 1 3261 FA1S $T=572880 457080 0 180 $X=561100 $Y=451660
X4048 3381 2 3358 3347 3415 1 3400 FA1S $T=564820 477240 1 0 $X=564820 $Y=471820
X4049 3390 2 406 3416 421 1 3419 FA1S $T=566680 537720 1 0 $X=566680 $Y=532300
X4050 3406 2 3425 3391 3432 1 3380 FA1S $T=581560 457080 1 180 $X=569780 $Y=456700
X4051 3409 2 3423 3401 3383 1 3461 FA1S $T=572260 497400 0 0 $X=572260 $Y=497020
X4052 3433 2 438 425 3377 1 3468 FA1S $T=573500 527640 1 0 $X=573500 $Y=522220
X4053 3446 2 3411 428 3434 1 3491 FA1S $T=576600 507480 0 0 $X=576600 $Y=507100
X4054 3451 2 3436 3419 3446 1 3482 FA1S $T=577220 517560 1 0 $X=577220 $Y=512140
X4055 3474 2 3503 3494 3486 1 3435 FA1S $T=590240 467160 0 180 $X=578460 $Y=461740
X4056 3457 2 3490 3440 3407 1 3486 FA1S $T=578460 477240 0 0 $X=578460 $Y=476860
X4057 3475 2 436 3499 432 1 3436 FA1S $T=590240 537720 0 180 $X=578460 $Y=532300
X4058 3489 2 3448 3457 3508 1 3439 FA1S $T=592720 477240 0 180 $X=580940 $Y=471820
X4059 3504 2 3480 3467 3396 1 3508 FA1S $T=585900 497400 1 0 $X=585900 $Y=491980
X4060 3517 2 3546 3504 3491 1 3552 FA1S $T=587140 487320 0 0 $X=587140 $Y=486940
X4061 3523 2 3514 3555 3575 1 3560 FA1S $T=589000 376440 1 0 $X=589000 $Y=371020
X4062 3546 2 3553 3577 3531 1 3481 FA1S $T=602020 477240 1 180 $X=590240 $Y=476860
X4063 457 2 439 3454 3559 1 3514 FA1S $T=602640 366360 1 180 $X=590860 $Y=365980
X4064 456 2 455 3475 3390 1 3534 FA1S $T=592720 537720 1 0 $X=592720 $Y=532300
X4065 3582 2 3463 3459 3661 1 3649 FA1S $T=598300 376440 0 0 $X=598300 $Y=376060
X4066 3565 2 3582 3571 3618 1 3593 FA1S $T=598300 386520 0 0 $X=598300 $Y=386140
X4067 3598 2 3104 3629 3604 1 3684 FA1S $T=600160 447000 0 0 $X=600160 $Y=446620
X4068 3575 2 3591 3683 3633 1 3571 FA1S $T=613800 376440 0 180 $X=602020 $Y=371020
X4069 3607 2 3605 3020 3596 1 3655 FA1S $T=602020 467160 0 0 $X=602020 $Y=466780
X4070 3612 2 3645 3644 3597 1 3670 FA1S $T=602640 416760 1 0 $X=602640 $Y=411340
X4071 3634 2 3592 3662 3652 1 3597 FA1S $T=616280 396600 0 180 $X=604500 $Y=391180
X4072 3627 2 407 3594 3616 1 3679 FA1S $T=604500 497400 0 0 $X=604500 $Y=497020
X4073 3583 2 3634 3611 3612 1 3635 FA1S $T=605740 396600 0 0 $X=605740 $Y=396220
X4074 3638 2 3615 3622 3609 1 3701 FA1S $T=606360 477240 0 0 $X=606360 $Y=476860
X4075 3647 2 3648 3632 3628 1 3697 FA1S $T=607600 537720 1 0 $X=607600 $Y=532300
X4076 3645 2 3493 3464 3708 1 3712 FA1S $T=609460 406680 1 0 $X=609460 $Y=401260
X4077 3618 2 3720 3649 3711 1 3611 FA1S $T=623720 386520 0 180 $X=611940 $Y=381100
X4078 3673 2 3676 3674 3607 1 3716 FA1S $T=613800 457080 1 0 $X=613800 $Y=451660
X4079 3721 2 3756 3712 3714 1 3681 FA1S $T=628060 416760 0 180 $X=616280 $Y=411340
X4080 3710 2 3646 3677 3746 1 3753 FA1S $T=616280 517560 1 0 $X=616280 $Y=512140
X4081 3642 2 3721 3670 3743 1 3664 FA1S $T=628680 416760 1 180 $X=616900 $Y=416380
X4082 3678 2 3681 3752 3722 1 3692 FA1S $T=629920 426840 0 180 $X=618140 $Y=421420
X4083 3724 2 3689 3700 3653 1 3769 FA1S $T=618760 477240 1 0 $X=618760 $Y=471820
X4084 3725 2 3704 3627 3701 1 3783 FA1S $T=618760 487320 1 0 $X=618760 $Y=481900
X4085 3726 2 3679 3705 3710 1 3781 FA1S $T=618760 497400 1 0 $X=618760 $Y=491980
X4086 3727 2 3663 3640 470 1 3763 FA1S $T=618760 527640 0 0 $X=618760 $Y=527260
X4087 3705 2 3702 3643 3637 1 3764 FA1S $T=619380 507480 1 0 $X=619380 $Y=502060
X4088 3740 2 3697 476 3763 1 481 FA1S $T=620620 537720 1 0 $X=620620 $Y=532300
X4089 3717 2 3685 3688 3732 1 3786 FA1S $T=621240 467160 0 0 $X=621240 $Y=466780
X4090 3747 2 3764 3647 3753 1 3785 FA1S $T=622480 507480 0 0 $X=622480 $Y=507100
X4091 3749 2 3691 3639 3682 1 3787 FA1S $T=623100 487320 0 0 $X=623100 $Y=486940
X4092 3767 2 3738 3779 3814 1 3802 FA1S $T=627440 406680 0 0 $X=627440 $Y=406300
X4093 3743 2 3767 3816 3810 1 3752 FA1S $T=641700 416760 0 180 $X=629920 $Y=411340
X4094 3810 2 3806 3827 3802 1 3768 FA1S $T=643560 416760 1 180 $X=631780 $Y=416380
X4095 3806 2 3421 3420 3792 1 3845 FA1S $T=633020 426840 1 0 $X=633020 $Y=421420
X4096 3722 2 3862 3896 3768 1 3803 FA1S $T=648520 426840 1 180 $X=636740 $Y=426460
X4097 3723 2 3882 3803 3848 1 3772 FA1S $T=648520 436920 0 180 $X=636740 $Y=431500
X4098 3856 2 3855 3822 3846 1 3901 FA1S $T=642320 416760 1 0 $X=642320 $Y=411340
X4099 3885 2 3570 3443 3812 1 3937 FA1S $T=646040 416760 0 0 $X=646040 $Y=416380
X4100 3896 2 3861 3845 3903 1 3939 FA1S $T=648520 426840 1 0 $X=648520 $Y=421420
X4101 3905 2 3891 3808 3868 1 3949 FA1S $T=649760 376440 0 0 $X=649760 $Y=376060
X4102 3848 2 3939 3938 3892 1 3969 FA1S $T=650380 436920 0 0 $X=650380 $Y=436540
X4103 3882 2 3946 3856 3940 1 3892 FA1S $T=663400 436920 0 180 $X=651620 $Y=431500
X4104 3938 2 3885 3968 3978 1 4014 FA1S $T=660300 416760 0 0 $X=660300 $Y=416380
X4105 3793 2 4024 3969 4000 1 3745 FA1S $T=675800 436920 1 180 $X=664020 $Y=436540
X4106 4009 2 3975 3905 4032 1 4061 FA1S $T=669600 376440 0 0 $X=669600 $Y=376060
X4107 4000 2 4014 4009 4074 1 4025 FA1S $T=673940 416760 1 0 $X=673940 $Y=411340
X4108 4024 2 4010 3901 4076 1 4074 FA1S $T=675180 406680 0 0 $X=675180 $Y=406300
X4109 4051 2 543 540 542 1 551 FA1S $T=675800 366360 0 0 $X=675800 $Y=365980
X4110 4008 2 527 4026 4051 1 4093 FA1S $T=677660 386520 1 0 $X=677660 $Y=381100
X4111 4092 2 4043 3949 4059 1 562 FA1S $T=686960 376440 1 0 $X=686960 $Y=371020
X4112 1206 17 1211 2 1 XNR2HS $T=225680 406680 0 180 $X=220100 $Y=401260
X4113 1208 1207 1213 2 1 XNR2HS $T=225680 457080 1 180 $X=220100 $Y=456700
X4114 1217 1219 1214 2 1 XNR2HS $T=225680 497400 1 180 $X=220100 $Y=497020
X4115 11 15 1236 2 1 XNR2HS $T=221960 376440 1 0 $X=221960 $Y=371020
X4116 1208 17 1229 2 1 XNR2HS $T=228780 457080 0 180 $X=223200 $Y=451660
X4117 1206 15 1244 2 1 XNR2HS $T=223820 406680 0 0 $X=223820 $Y=406300
X4118 7 1207 1245 2 1 XNR2HS $T=223820 447000 0 0 $X=223820 $Y=446620
X4119 1205 21 1247 2 1 XNR2HS $T=224440 376440 0 0 $X=224440 $Y=376060
X4120 1230 15 1249 2 1 XNR2HS $T=225060 447000 1 0 $X=225060 $Y=441580
X4121 1206 1207 1253 2 1 XNR2HS $T=225680 416760 0 0 $X=225680 $Y=416380
X4122 1230 24 1254 2 1 XNR2HS $T=225680 426840 1 0 $X=225680 $Y=421420
X4123 1206 24 1252 2 1 XNR2HS $T=226300 386520 0 0 $X=226300 $Y=386140
X4124 1230 17 1257 2 1 XNR2HS $T=226300 436920 1 0 $X=226300 $Y=431500
X4125 1208 15 1258 2 1 XNR2HS $T=226300 457080 0 0 $X=226300 $Y=456700
X4126 1217 1250 1265 2 1 XNR2HS $T=227540 497400 1 0 $X=227540 $Y=491980
X4127 25 1243 1277 2 1 XNR2HS $T=230640 497400 0 0 $X=230640 $Y=497020
X4128 1230 32 1276 2 1 XNR2HS $T=237460 416760 1 180 $X=231880 $Y=416380
X4129 1217 24 1290 2 1 XNR2HS $T=231880 477240 0 0 $X=231880 $Y=476860
X4130 1269 24 1295 2 1 XNR2HS $T=232500 447000 1 0 $X=232500 $Y=441580
X4131 1264 32 1283 2 1 XNR2HS $T=238700 477240 0 180 $X=233120 $Y=471820
X4132 1269 32 1313 2 1 XNR2HS $T=236220 436920 0 0 $X=236220 $Y=436540
X4133 1328 1323 1306 2 1 XNR2HS $T=243040 416760 0 180 $X=237460 $Y=411340
X4134 1269 35 1325 2 1 XNR2HS $T=238080 447000 1 0 $X=238080 $Y=441580
X4135 1264 35 1307 2 1 XNR2HS $T=238080 477240 0 0 $X=238080 $Y=476860
X4136 1305 1250 1327 2 1 XNR2HS $T=238080 507480 0 0 $X=238080 $Y=507100
X4137 1338 32 1317 2 1 XNR2HS $T=244900 497400 1 180 $X=239320 $Y=497020
X4138 1343 32 1282 2 1 XNR2HS $T=246140 386520 0 180 $X=240560 $Y=381100
X4139 1305 1243 1351 2 1 XNR2HS $T=242420 517560 1 0 $X=242420 $Y=512140
X4140 1264 46 1341 2 1 XNR2HS $T=250480 467160 0 180 $X=244900 $Y=461740
X4141 1338 41 1361 2 1 XNR2HS $T=244900 487320 1 0 $X=244900 $Y=481900
X4142 1343 35 1302 2 1 XNR2HS $T=246140 386520 1 0 $X=246140 $Y=381100
X4143 1353 35 1291 2 1 XNR2HS $T=246140 406680 0 0 $X=246140 $Y=406300
X4144 1338 35 1365 2 1 XNR2HS $T=246140 497400 1 0 $X=246140 $Y=491980
X4145 1348 48 1308 2 1 XNR2HS $T=252340 426840 0 180 $X=246760 $Y=421420
X4146 1338 46 1367 2 1 XNR2HS $T=246760 477240 0 0 $X=246760 $Y=476860
X4147 1353 46 1363 2 1 XNR2HS $T=253580 396600 1 180 $X=248000 $Y=396220
X4148 1264 41 1345 2 1 XNR2HS $T=248000 467160 0 0 $X=248000 $Y=466780
X4149 1338 48 1371 2 1 XNR2HS $T=248000 477240 1 0 $X=248000 $Y=471820
X4150 1359 38 1372 2 1 XNR2HS $T=248000 507480 1 0 $X=248000 $Y=502060
X4151 1301 1366 53 2 1 XNR2HS $T=248620 386520 0 0 $X=248620 $Y=386140
X4152 1348 46 1337 2 1 XNR2HS $T=254200 426840 1 180 $X=248620 $Y=426460
X4153 1305 1319 1375 2 1 XNR2HS $T=248620 517560 1 0 $X=248620 $Y=512140
X4154 1348 41 1360 2 1 XNR2HS $T=251100 436920 1 0 $X=251100 $Y=431500
X4155 1264 48 1326 2 1 XNR2HS $T=251100 457080 0 0 $X=251100 $Y=456700
X4156 1343 41 1389 2 1 XNR2HS $T=251720 376440 0 0 $X=251720 $Y=376060
X4157 1353 41 1368 2 1 XNR2HS $T=259160 406680 0 180 $X=253580 $Y=401260
X4158 1353 48 1378 2 1 XNR2HS $T=259780 396600 1 180 $X=254200 $Y=396220
X4159 1390 1355 1412 2 1 XNR2HS $T=256680 457080 0 0 $X=256680 $Y=456700
X4160 56 47 57 2 1 XNR2HS $T=256680 537720 1 0 $X=256680 $Y=532300
X4161 1343 46 1421 2 1 XNR2HS $T=257920 376440 1 0 $X=257920 $Y=371020
X4162 1431 1408 1415 2 1 XNR2HS $T=264740 477240 0 180 $X=259160 $Y=471820
X4163 1420 50 1432 2 1 XNR2HS $T=260400 517560 1 0 $X=260400 $Y=512140
X4164 1420 60 1434 2 1 XNR2HS $T=261020 497400 1 0 $X=261020 $Y=491980
X4165 1420 43 1435 2 1 XNR2HS $T=261020 507480 1 0 $X=261020 $Y=502060
X4166 1397 1405 62 2 1 XNR2HS $T=261640 366360 0 0 $X=261640 $Y=365980
X4167 1420 1386 1442 2 1 XNR2HS $T=262260 507480 0 0 $X=262260 $Y=507100
X4168 56 38 1444 2 1 XNR2HS $T=262880 527640 1 0 $X=262880 $Y=522220
X4169 56 39 1445 2 1 XNR2HS $T=262880 537720 1 0 $X=262880 $Y=532300
X4170 1413 48 1436 2 1 XNR2HS $T=267840 386520 1 0 $X=267840 $Y=381100
X4171 1472 1469 1455 2 1 XNR2HS $T=273420 477240 1 180 $X=267840 $Y=476860
X4172 1420 64 1462 2 1 XNR2HS $T=271560 497400 0 0 $X=271560 $Y=497020
X4173 70 60 1488 2 1 XNR2HS $T=272800 517560 0 0 $X=272800 $Y=517180
X4174 76 1522 1506 2 1 XNR2HS $T=283960 507480 1 180 $X=278380 $Y=507100
X4175 70 39 75 2 1 XNR2HS $T=278380 537720 1 0 $X=278380 $Y=532300
X4176 70 64 1523 2 1 XNR2HS $T=279620 527640 1 0 $X=279620 $Y=522220
X4177 1691 1722 1760 2 1 XNR2HS $T=312480 406680 1 0 $X=312480 $Y=401260
X4178 1730 1677 1763 2 1 XNR2HS $T=312480 457080 1 0 $X=312480 $Y=451660
X4179 110 109 1741 2 1 XNR2HS $T=318680 537720 0 180 $X=313100 $Y=532300
X4180 1729 1765 1773 2 1 XNR2HS $T=314960 416760 0 0 $X=314960 $Y=416380
X4181 1767 1749 1777 2 1 XNR2HS $T=315580 477240 0 0 $X=315580 $Y=476860
X4182 1752 1709 1811 2 1 XNR2HS $T=321160 396600 0 0 $X=321160 $Y=396220
X4183 1783 1817 1843 2 1 XNR2HS $T=326740 487320 0 0 $X=326740 $Y=486940
X4184 2049 2019 2073 2 1 XNR2HS $T=365800 497400 0 0 $X=365800 $Y=497020
X4185 2220 2224 2239 2 1 XNR2HS $T=391220 497400 0 0 $X=391220 $Y=497020
X4186 2372 227 2407 2 1 XNR2HS $T=429660 416760 0 180 $X=424080 $Y=411340
X4187 232 227 2424 2 1 XNR2HS $T=435240 376440 0 180 $X=429660 $Y=371020
X4188 234 227 2443 2 1 XNR2HS $T=435240 386520 1 180 $X=429660 $Y=386140
X4189 235 227 2432 2 1 XNR2HS $T=435240 406680 0 180 $X=429660 $Y=401260
X4190 2446 2423 2461 2 1 XNR2HS $T=431520 487320 0 0 $X=431520 $Y=486940
X4191 2477 2480 2491 2 1 XNR2HS $T=435860 507480 1 0 $X=435860 $Y=502060
X4192 2505 2499 2415 2 1 XNR2HS $T=442060 447000 1 180 $X=436480 $Y=446620
X4193 235 242 2496 2 1 XNR2HS $T=437100 376440 0 0 $X=437100 $Y=376060
X4194 246 242 2525 2 1 XNR2HS $T=440200 406680 1 0 $X=440200 $Y=401260
X4195 2521 2535 2520 2 1 XNR2HS $T=447640 447000 1 180 $X=442060 $Y=446620
X4196 2499 2542 2535 2 1 XNR2HS $T=445160 457080 1 0 $X=445160 $Y=451660
X4197 245 2528 2543 2 1 XNR2HS $T=445160 527640 0 0 $X=445160 $Y=527260
X4198 2380 2576 2565 2 1 XNR2HS $T=455080 386520 0 180 $X=449500 $Y=381100
X4199 2380 242 2539 2 1 XNR2HS $T=456320 406680 0 180 $X=450740 $Y=401260
X4200 264 242 2552 2 1 XNR2HS $T=456940 366360 1 180 $X=451360 $Y=365980
X4201 2568 2579 2589 2 1 XNR2HS $T=451980 436920 1 0 $X=451980 $Y=431500
X4202 2560 2569 2573 2 1 XNR2HS $T=451980 436920 0 0 $X=451980 $Y=436540
X4203 2574 242 2540 2 1 XNR2HS $T=458180 416760 0 180 $X=452600 $Y=411340
X4204 2575 2594 2569 2 1 XNR2HS $T=458180 447000 1 180 $X=452600 $Y=446620
X4205 246 2576 2599 2 1 XNR2HS $T=453840 396600 1 0 $X=453840 $Y=391180
X4206 2601 2610 2579 2 1 XNR2HS $T=460660 447000 0 180 $X=455080 $Y=441580
X4207 264 257 267 2 1 XNR2HS $T=466240 366360 1 180 $X=460660 $Y=365980
X4208 2665 2658 2616 2 1 XNR2HS $T=468720 447000 0 180 $X=463140 $Y=441580
X4209 284 2576 2641 2 1 XNR2HS $T=471820 386520 1 180 $X=466240 $Y=386140
X4210 2657 2673 2685 2 1 XNR2HS $T=466860 436920 1 0 $X=466860 $Y=431500
X4211 284 272 280 2 1 XNR2HS $T=473060 366360 1 180 $X=467480 $Y=365980
X4212 2690 2688 2673 2 1 XNR2HS $T=470580 436920 0 0 $X=470580 $Y=436540
X4213 2764 2769 2773 2 1 XNR2HS $T=482980 436920 0 0 $X=482980 $Y=436540
X4214 3202 3195 2769 2 1 XNR2HS $T=541880 436920 1 180 $X=536300 $Y=436540
X4215 3220 3203 2674 2 1 XNR2HS $T=544980 447000 1 180 $X=539400 $Y=446620
X4216 3328 3325 3229 2 1 XNR2HS $T=561720 447000 0 180 $X=556140 $Y=441580
X4217 3352 3351 3319 2 1 XNR2HS $T=566060 436920 1 180 $X=560480 $Y=436540
X4218 3405 3402 3331 2 1 XNR2HS $T=575360 376440 1 180 $X=569780 $Y=376060
X4219 3453 3450 3382 2 1 XNR2HS $T=583420 447000 0 180 $X=577840 $Y=441580
X4220 3455 3438 3321 2 1 XNR2HS $T=584040 396600 1 180 $X=578460 $Y=396220
X4221 3460 3456 3444 2 1 XNR2HS $T=584660 436920 1 180 $X=579080 $Y=436540
X4222 3469 3465 3392 2 1 XNR2HS $T=585900 416760 1 180 $X=580320 $Y=416380
X4223 3449 3444 443 2 1 XNR2HS $T=580940 426840 0 0 $X=580940 $Y=426460
X4224 3477 3472 3387 2 1 XNR2HS $T=587140 416760 0 180 $X=581560 $Y=411340
X4225 3496 3487 3327 2 1 XNR2HS $T=589620 396600 0 180 $X=584040 $Y=391180
X4226 3497 3483 3356 2 1 XNR2HS $T=589620 396600 1 180 $X=584040 $Y=396220
X4227 3498 3488 3385 2 1 XNR2HS $T=589620 426840 0 180 $X=584040 $Y=421420
X4228 3516 3515 3336 2 1 XNR2HS $T=592720 426840 1 180 $X=587140 $Y=426460
X4229 3562 3458 3506 2 1 XNR2HS $T=603880 497400 0 180 $X=598300 $Y=491980
X4230 3561 3574 3585 2 1 XNR2HS $T=599540 507480 0 0 $X=599540 $Y=507100
X4231 3556 3578 3589 2 1 XNR2HS $T=600160 447000 1 0 $X=600160 $Y=441580
X4232 3603 3599 3363 2 1 XNR2HS $T=606980 426840 0 180 $X=601400 $Y=421420
X4233 3589 3600 3581 2 1 XNR2HS $T=606980 436920 1 180 $X=601400 $Y=436540
X4234 3554 3585 466 2 1 XNR2HS $T=606980 436920 0 0 $X=606980 $Y=436540
X4235 3620 3598 3651 2 1 XNR2HS $T=608840 447000 1 0 $X=608840 $Y=441580
X4236 468 467 3625 2 1 XNR2HS $T=615040 366360 1 180 $X=609460 $Y=365980
X4237 2664 467 3660 2 1 XNR2HS $T=610700 386520 0 0 $X=610700 $Y=386140
X4238 2966 467 3698 2 1 XNR2HS $T=616900 386520 0 0 $X=616900 $Y=386140
X4239 3651 3669 3709 2 1 XNR2HS $T=616900 436920 1 0 $X=616900 $Y=431500
X4240 131 467 3687 2 1 XNR2HS $T=624960 366360 1 180 $X=619380 $Y=365980
X4241 472 3709 3713 2 1 XNR2HS $T=628060 396600 0 180 $X=622480 $Y=391180
X4242 2399 3709 3751 2 1 XNR2HS $T=624340 396600 0 0 $X=624340 $Y=396220
X4243 475 474 3719 2 1 XNR2HS $T=630540 366360 1 180 $X=624960 $Y=365980
X4244 3716 3699 3762 2 1 XNR2HS $T=626200 457080 1 0 $X=626200 $Y=451660
X4245 3610 480 3601 2 1 XNR2HS $T=633640 517560 1 180 $X=628060 $Y=517180
X4246 482 3775 3750 2 1 XNR2HS $T=634260 376440 1 180 $X=628680 $Y=376060
X4247 483 3776 3744 2 1 XNR2HS $T=634260 386520 0 180 $X=628680 $Y=381100
X4248 225 3760 3774 2 1 XNR2HS $T=628680 396600 1 0 $X=628680 $Y=391180
X4249 3777 3773 3761 2 1 XNR2HS $T=634260 447000 0 180 $X=628680 $Y=441580
X4250 468 3775 3729 2 1 XNR2HS $T=634880 376440 0 180 $X=629300 $Y=371020
X4251 3755 3718 3777 2 1 XNR2HS $T=629300 447000 0 0 $X=629300 $Y=446620
X4252 2664 3776 3782 2 1 XNR2HS $T=639840 386520 1 180 $X=634260 $Y=386140
X4253 3715 3798 3807 2 1 XNR2HS $T=634260 507480 0 0 $X=634260 $Y=507100
X4254 225 3776 3813 2 1 XNR2HS $T=635500 386520 1 0 $X=635500 $Y=381100
X4255 3799 3805 3798 2 1 XNR2HS $T=636120 517560 0 0 $X=636120 $Y=517180
X4256 2399 3776 3826 2 1 XNR2HS $T=637980 396600 1 0 $X=637980 $Y=391180
X4257 493 3796 3821 2 1 XNR2HS $T=639840 376440 1 0 $X=639840 $Y=371020
X4258 493 3775 495 2 1 XNR2HS $T=641700 366360 0 0 $X=641700 $Y=365980
X4259 499 496 3832 2 1 XNR2HS $T=647280 537720 0 180 $X=641700 $Y=532300
X4260 2966 3776 3836 2 1 XNR2HS $T=642940 406680 1 0 $X=642940 $Y=401260
X4261 472 3776 3858 2 1 XNR2HS $T=643560 396600 1 0 $X=643560 $Y=391180
X4262 3832 3819 3859 2 1 XNR2HS $T=643560 517560 0 0 $X=643560 $Y=517180
X4263 3850 3828 3864 2 1 XNR2HS $T=644180 447000 0 0 $X=644180 $Y=446620
X4264 3847 3852 3866 2 1 XNR2HS $T=644180 477240 0 0 $X=644180 $Y=476860
X4265 3835 3817 3887 2 1 XNR2HS $T=647280 457080 1 0 $X=647280 $Y=451660
X4266 3870 3871 3889 2 1 XNR2HS $T=647280 507480 1 0 $X=647280 $Y=502060
X4267 482 3894 3875 2 1 XNR2HS $T=654100 386520 0 180 $X=648520 $Y=381100
X4268 3864 3879 3877 2 1 XNR2HS $T=648520 447000 1 0 $X=648520 $Y=441580
X4269 3902 3878 3884 2 1 XNR2HS $T=654720 527640 0 180 $X=649140 $Y=522220
X4270 475 3894 3876 2 1 XNR2HS $T=655340 396600 0 180 $X=649760 $Y=391180
X4271 501 3766 3900 2 1 XNR2HS $T=650380 517560 1 0 $X=650380 $Y=512140
X4272 3884 3834 3909 2 1 XNR2HS $T=651000 517560 0 0 $X=651000 $Y=517180
X4273 3887 3880 509 2 1 XNR2HS $T=652240 447000 0 0 $X=652240 $Y=446620
X4274 3900 506 510 2 1 XNR2HS $T=652860 507480 1 0 $X=652860 $Y=502060
X4275 514 509 3908 2 1 XNR2HS $T=659060 406680 0 180 $X=653480 $Y=401260
X4276 3889 3911 3922 2 1 XNR2HS $T=653480 497400 0 0 $X=653480 $Y=497020
X4277 482 508 3929 2 1 XNR2HS $T=654100 386520 1 0 $X=654100 $Y=381100
X4278 3890 3898 3923 2 1 XNR2HS $T=654720 477240 0 0 $X=654720 $Y=476860
X4279 482 511 3933 2 1 XNR2HS $T=655340 376440 1 0 $X=655340 $Y=371020
X4280 3923 3910 3934 2 1 XNR2HS $T=655340 467160 0 0 $X=655340 $Y=466780
X4281 475 508 3914 2 1 XNR2HS $T=663400 386520 1 180 $X=657820 $Y=386140
X4282 483 509 3931 2 1 XNR2HS $T=664640 406680 0 180 $X=659060 $Y=401260
X4283 472 508 524 2 1 XNR2HS $T=662780 366360 0 0 $X=662780 $Y=365980
X4284 483 3894 3976 2 1 XNR2HS $T=662780 396600 0 0 $X=662780 $Y=396220
X4285 475 510 3977 2 1 XNR2HS $T=662780 426840 0 0 $X=662780 $Y=426460
X4286 2966 508 3959 2 1 XNR2HS $T=668980 386520 1 180 $X=663400 $Y=386140
X4287 514 3894 3915 2 1 XNR2HS $T=664020 396600 1 0 $X=664020 $Y=391180
X4288 2664 509 3950 2 1 XNR2HS $T=671460 406680 1 180 $X=665880 $Y=406300
X4289 514 511 3994 2 1 XNR2HS $T=667740 376440 1 0 $X=667740 $Y=371020
X4290 2664 3894 3997 2 1 XNR2HS $T=668360 396600 0 0 $X=668360 $Y=396220
X4291 483 511 532 2 1 XNR2HS $T=668980 366360 0 0 $X=668980 $Y=365980
X4292 2966 3894 533 2 1 XNR2HS $T=668980 386520 0 0 $X=668980 $Y=386140
X4293 2667 2721 2771 1 2 2847 OA12 $T=492900 487320 1 0 $X=492900 $Y=481900
X4294 2901 339 2935 1 2 2973 OA12 $T=510260 416760 1 0 $X=510260 $Y=411340
X4295 3410 422 3397 1 2 3297 OA12 $T=575360 386520 0 180 $X=571640 $Y=381100
X4296 3437 3431 3427 1 2 3397 OA12 $T=579700 376440 1 180 $X=575980 $Y=376060
X4297 3426 3442 427 1 2 3427 OA12 $T=582180 376440 0 180 $X=578460 $Y=371020
X4298 1235 1 1211 1222 1251 1244 2 OAI22S $T=226300 406680 1 0 $X=226300 $Y=401260
X4299 1235 1 1252 1222 1248 1211 2 OAI22S $T=231260 396600 0 180 $X=227540 $Y=391180
X4300 26 1 27 28 1272 1236 2 OAI22S $T=230020 366360 0 0 $X=230020 $Y=365980
X4301 1235 1 1244 1222 1263 1253 2 OAI22S $T=233740 406680 1 180 $X=230020 $Y=406300
X4302 26 1 1236 1226 1266 1247 2 OAI22S $T=234360 376440 0 180 $X=230640 $Y=371020
X4303 1280 1 1276 1221 1260 1254 2 OAI22S $T=234980 426840 0 180 $X=231260 $Y=421420
X4304 1280 1 1254 1221 1273 1257 2 OAI22S $T=235600 426840 1 180 $X=231880 $Y=426460
X4305 1280 1 1257 1221 1274 1249 2 OAI22S $T=235600 436920 1 180 $X=231880 $Y=436540
X4306 1280 1 1249 1221 1275 1245 2 OAI22S $T=235600 447000 1 180 $X=231880 $Y=446620
X4307 1241 1 1258 1240 1271 1213 2 OAI22S $T=235600 467160 0 180 $X=231880 $Y=461740
X4308 1235 1 1282 1222 1279 1252 2 OAI22S $T=236220 386520 0 180 $X=232500 $Y=381100
X4309 1293 1 1265 1278 1281 1277 2 OAI22S $T=236840 487320 1 180 $X=233120 $Y=486940
X4310 1280 1 1291 1221 1285 1276 2 OAI22S $T=237460 406680 1 180 $X=233740 $Y=406300
X4311 1262 1 1294 1299 1301 1308 2 OAI22S $T=234980 426840 1 0 $X=234980 $Y=421420
X4312 1293 1 1277 1296 1292 1214 2 OAI22S $T=238700 497400 0 180 $X=234980 $Y=491980
X4313 1235 1 1302 1222 33 1282 2 OAI22S $T=239940 386520 0 180 $X=236220 $Y=381100
X4314 1241 1 1229 1240 1311 1258 2 OAI22S $T=236220 467160 1 0 $X=236220 $Y=461740
X4315 1314 1 1307 1297 1303 1283 2 OAI22S $T=240560 467160 1 180 $X=236840 $Y=466780
X4316 1294 1 1313 1240 1310 1295 2 OAI22S $T=241800 436920 0 180 $X=238080 $Y=431500
X4317 1294 1 1308 1299 1329 1337 2 OAI22S $T=239320 426840 1 0 $X=239320 $Y=421420
X4318 1314 1 1283 1278 1330 1290 2 OAI22S $T=239320 477240 1 0 $X=239320 $Y=471820
X4319 1309 1 1295 1240 1318 1229 2 OAI22S $T=243660 447000 1 180 $X=239940 $Y=446620
X4320 1316 1 1320 1297 1328 1326 2 OAI22S $T=239940 457080 0 0 $X=239940 $Y=456700
X4321 1320 1 1326 1297 1335 1341 2 OAI22S $T=240560 467160 1 0 $X=240560 $Y=461740
X4322 1314 1 1290 1278 1324 1265 2 OAI22S $T=244280 487320 0 180 $X=240560 $Y=481900
X4323 1316 1 1278 1286 1333 1314 2 OAI22S $T=245520 487320 1 180 $X=241800 $Y=486940
X4324 1309 1 1325 1299 1334 1313 2 OAI22S $T=246140 436920 0 180 $X=242420 $Y=431500
X4325 1314 1 1345 1278 1342 1307 2 OAI22S $T=247380 477240 0 180 $X=243660 $Y=471820
X4326 1309 1 1337 1299 1323 1360 2 OAI22S $T=244280 426840 0 0 $X=244280 $Y=426460
X4327 1262 1 1240 1349 1350 1309 2 OAI22S $T=244280 447000 0 0 $X=244280 $Y=446620
X4328 1320 1 1341 1297 1355 1345 2 OAI22S $T=244280 467160 0 0 $X=244280 $Y=466780
X4329 1309 1 1360 1299 1357 1325 2 OAI22S $T=250480 436920 0 180 $X=246760 $Y=431500
X4330 1322 1 1363 1346 1366 1368 2 OAI22S $T=247380 396600 1 0 $X=247380 $Y=391180
X4331 1322 1 1378 1346 54 1363 2 OAI22S $T=255440 396600 0 180 $X=251720 $Y=391180
X4332 1322 1 1368 1346 1379 1291 2 OAI22S $T=256060 406680 1 180 $X=252340 $Y=406300
X4333 1370 1 1365 1384 1373 1317 2 OAI22S $T=252340 487320 0 0 $X=252340 $Y=486940
X4334 1370 1 1361 1384 1381 1365 2 OAI22S $T=256680 477240 1 180 $X=252960 $Y=476860
X4335 1396 1 1370 1384 1390 1371 2 OAI22S $T=257920 467160 0 180 $X=254200 $Y=461740
X4336 1385 1 1351 1392 1393 1375 2 OAI22S $T=257920 517560 1 180 $X=254200 $Y=517180
X4337 1370 1 1371 1384 1398 1367 2 OAI22S $T=254820 477240 1 0 $X=254820 $Y=471820
X4338 1385 1 1317 1392 1399 1372 2 OAI22S $T=254820 497400 0 0 $X=254820 $Y=497020
X4339 1385 1 1327 1392 1391 1351 2 OAI22S $T=258540 507480 1 180 $X=254820 $Y=507100
X4340 1414 1 1322 1346 1397 1378 2 OAI22S $T=259780 396600 0 180 $X=256060 $Y=391180
X4341 1394 1 1389 1289 1401 1302 2 OAI22S $T=261020 376440 1 180 $X=257300 $Y=376060
X4342 1385 1 1372 1392 1404 1327 2 OAI22S $T=261020 507480 0 180 $X=257300 $Y=502060
X4343 1370 1 1367 1384 1408 1361 2 OAI22S $T=261640 477240 1 180 $X=257920 $Y=476860
X4344 1396 1 1392 1387 1419 1385 2 OAI22S $T=258540 507480 0 0 $X=258540 $Y=507100
X4345 1414 1 1346 1417 1424 1322 2 OAI22S $T=260400 406680 0 0 $X=260400 $Y=406300
X4346 1394 1 1421 1289 1405 1389 2 OAI22S $T=265360 376440 1 180 $X=261640 $Y=376060
X4347 1433 1 1289 1428 1423 1394 2 OAI22S $T=265980 386520 0 180 $X=262260 $Y=381100
X4348 1394 1 1436 1289 61 1421 2 OAI22S $T=267220 376440 0 180 $X=263500 $Y=371020
X4349 1446 1 1434 1453 1449 1462 2 OAI22S $T=266600 487320 0 0 $X=266600 $Y=486940
X4350 63 1 1432 65 1456 1444 2 OAI22S $T=266600 517560 1 0 $X=266600 $Y=512140
X4351 1433 1 1394 1289 66 1436 2 OAI22S $T=267220 376440 1 0 $X=267220 $Y=371020
X4352 1458 1 1446 1453 1431 1434 2 OAI22S $T=270940 487320 0 180 $X=267220 $Y=481900
X4353 1446 1 1435 1453 1450 1442 2 OAI22S $T=270940 497400 1 180 $X=267220 $Y=497020
X4354 1446 1 1442 1453 1451 1432 2 OAI22S $T=270940 507480 0 180 $X=267220 $Y=502060
X4355 63 1 1444 65 1463 1445 2 OAI22S $T=272800 527640 0 180 $X=269080 $Y=522220
X4356 1458 1 65 1457 1470 63 2 OAI22S $T=269080 527640 0 0 $X=269080 $Y=527260
X4357 63 1 1445 65 1464 57 2 OAI22S $T=272800 537720 0 180 $X=269080 $Y=532300
X4358 1446 1 1462 1453 1469 1435 2 OAI22S $T=274660 487320 1 180 $X=270940 $Y=486940
X4359 1481 1 1485 1486 1472 1488 2 OAI22S $T=274040 517560 1 0 $X=274040 $Y=512140
X4360 1481 1 1486 1493 1499 1485 2 OAI22S $T=275900 527640 0 0 $X=275900 $Y=527260
X4361 1485 1 1488 1486 1524 1523 2 OAI22S $T=282720 517560 1 0 $X=282720 $Y=512140
X4362 1485 1 1523 1486 1522 86 2 OAI22S $T=286440 517560 0 0 $X=286440 $Y=517180
X4363 85 1 83 80 1547 81 2 OAI22S $T=290780 537720 0 180 $X=287060 $Y=532300
X4364 79 1 90 1486 1574 88 2 OAI22S $T=295120 537720 0 180 $X=291400 $Y=532300
X4365 79 1 81 80 1597 75 2 OAI22S $T=299460 537720 0 180 $X=295740 $Y=532300
X4366 220 1 222 224 2419 2424 2 OAI22S $T=424700 366360 0 0 $X=424700 $Y=365980
X4367 226 1 2432 2415 2425 2407 2 OAI22S $T=430900 406680 1 180 $X=427180 $Y=406300
X4368 226 1 2424 224 2447 2443 2 OAI22S $T=429660 386520 1 0 $X=429660 $Y=381100
X4369 226 1 2443 224 2451 2432 2 OAI22S $T=430280 396600 0 0 $X=430280 $Y=396220
X4370 226 1 2407 2415 2455 2380 2 OAI22S $T=434000 416760 0 0 $X=434000 $Y=416380
X4371 2526 1 248 244 2502 2496 2 OAI22S $T=443920 366360 1 180 $X=440200 $Y=365980
X4372 2526 1 2525 2531 2509 2540 2 OAI22S $T=443300 416760 1 0 $X=443300 $Y=411340
X4373 2526 1 2552 2531 2524 2539 2 OAI22S $T=450120 396600 0 180 $X=446400 $Y=391180
X4374 2526 1 2539 2531 2548 2525 2 OAI22S $T=450120 406680 0 180 $X=446400 $Y=401260
X4375 2558 1 2529 2551 2550 2537 2 OAI22S $T=450120 426840 0 180 $X=446400 $Y=421420
X4376 2526 1 2496 244 2559 2552 2 OAI22S $T=447020 376440 0 0 $X=447020 $Y=376060
X4377 2586 1 193 2595 2578 2604 2 OAI22S $T=454460 487320 0 0 $X=454460 $Y=486940
X4378 2593 1 2565 2599 2602 262 2 OAI22S $T=455700 386520 0 0 $X=455700 $Y=386140
X4379 266 1 267 2565 2597 262 2 OAI22S $T=460660 366360 1 180 $X=456940 $Y=365980
X4380 2632 1 262 2622 2614 266 2 OAI22S $T=463140 396600 0 180 $X=459420 $Y=391180
X4381 2593 1 2599 2641 2639 262 2 OAI22S $T=466240 386520 0 180 $X=462520 $Y=381100
X4382 277 1 2656 2677 2681 273 2 OAI22S $T=466860 376440 0 0 $X=466860 $Y=376060
X4383 2485 1 289 2475 2694 2705 2 OAI22S $T=471200 406680 0 0 $X=471200 $Y=406300
X4384 2485 1 2025 2475 2718 2729 2 OAI22S $T=474920 416760 1 0 $X=474920 $Y=411340
X4385 3298 1 3327 3324 3311 3321 2 OAI22S $T=562340 406680 1 180 $X=558620 $Y=406300
X4386 2837 1 3297 3324 3337 3331 2 OAI22S $T=564820 416760 1 180 $X=561100 $Y=416380
X4387 3253 1 3297 3321 3339 3298 2 OAI22S $T=567920 416760 0 180 $X=564200 $Y=411340
X4388 3298 1 3365 3363 3342 2837 2 OAI22S $T=568540 426840 0 180 $X=564820 $Y=421420
X4389 3298 1 3336 3363 3369 3324 2 OAI22S $T=565440 416760 0 0 $X=565440 $Y=416380
X4390 3324 1 3336 3385 3348 3253 2 OAI22S $T=569160 426840 1 0 $X=569160 $Y=421420
X4391 2837 1 3321 3253 3389 3331 2 OAI22S $T=575360 416760 0 180 $X=571640 $Y=411340
X4392 3253 1 3392 2837 3384 3385 2 OAI22S $T=571640 416760 0 0 $X=571640 $Y=416380
X4393 459 1 460 461 3559 3625 2 OAI22S $T=605120 366360 0 0 $X=605120 $Y=365980
X4394 3625 1 460 461 3683 3687 2 OAI22S $T=615040 366360 0 0 $X=615040 $Y=365980
X4395 3687 1 460 3680 3661 3660 2 OAI22S $T=618760 376440 1 180 $X=615040 $Y=376060
X4396 3660 1 460 3680 3662 3698 2 OAI22S $T=616280 396600 1 0 $X=616280 $Y=391180
X4397 3698 1 3706 3680 3708 3713 2 OAI22S $T=618760 396600 0 0 $X=618760 $Y=396220
X4398 3729 1 3734 3728 3652 3744 2 OAI22S $T=623100 386520 0 0 $X=623100 $Y=386140
X4399 3750 1 3734 3728 3720 3729 2 OAI22S $T=628060 386520 0 180 $X=624340 $Y=381100
X4400 3719 1 3734 3728 3633 3750 2 OAI22S $T=624960 376440 1 0 $X=624960 $Y=371020
X4401 3744 1 3734 3728 3756 3782 2 OAI22S $T=629920 386520 0 0 $X=629920 $Y=386140
X4402 3713 1 3706 3754 3779 3774 2 OAI22S $T=630540 406680 1 0 $X=630540 $Y=401260
X4403 3774 1 485 3754 3792 3751 2 OAI22S $T=634260 396600 0 0 $X=634260 $Y=396220
X4404 490 1 485 489 3808 488 2 OAI22S $T=641080 366360 1 180 $X=637360 $Y=365980
X4405 3821 1 485 3754 3812 490 2 OAI22S $T=641700 376440 1 180 $X=637980 $Y=376060
X4406 3751 1 485 3754 3822 3821 2 OAI22S $T=638600 406680 1 0 $X=638600 $Y=401260
X4407 3782 1 3823 3831 3814 3836 2 OAI22S $T=639840 406680 0 0 $X=639840 $Y=406300
X4408 3813 1 498 497 3860 3826 2 OAI22S $T=644800 386520 1 0 $X=644800 $Y=381100
X4409 3836 1 3823 3831 3861 3858 2 OAI22S $T=644800 406680 0 0 $X=644800 $Y=406300
X4410 3826 1 498 497 3868 495 2 OAI22S $T=645420 376440 0 0 $X=645420 $Y=376060
X4411 3858 1 498 3831 3846 3813 2 OAI22S $T=649140 386520 1 180 $X=645420 $Y=386140
X4412 3873 1 3876 3881 3862 3875 2 OAI22S $T=648520 396600 0 0 $X=648520 $Y=396220
X4413 3873 1 3875 3881 3903 3915 2 OAI22S $T=652240 406680 0 0 $X=652240 $Y=406300
X4414 3908 1 3916 3921 3827 3931 2 OAI22S $T=654100 416760 1 0 $X=654100 $Y=411340
X4415 3914 1 512 3920 3644 3929 2 OAI22S $T=655960 396600 1 0 $X=655960 $Y=391180
X4416 3931 1 3916 3920 3946 3950 2 OAI22S $T=657820 416760 1 0 $X=657820 $Y=411340
X4417 3929 1 512 3920 3714 3908 2 OAI22S $T=662160 406680 1 180 $X=658440 $Y=406300
X4418 3950 1 512 3920 3968 3959 2 OAI22S $T=665880 406680 1 180 $X=662160 $Y=406300
X4419 3959 1 512 521 3975 524 2 OAI22S $T=664020 376440 0 0 $X=664020 $Y=376060
X4420 528 1 3977 525 3978 3933 2 OAI22S $T=670840 426840 0 180 $X=667120 $Y=421420
X4421 3917 1 3976 3881 4007 3997 2 OAI22S $T=670840 406680 1 0 $X=670840 $Y=401260
X4422 3917 1 3915 3881 4010 3976 2 OAI22S $T=671460 406680 0 0 $X=671460 $Y=406300
X4423 528 1 3933 539 4032 3994 2 OAI22S $T=674560 376440 1 0 $X=674560 $Y=371020
X4424 538 1 3997 3881 4043 533 2 OAI22S $T=677040 396600 0 0 $X=677040 $Y=396220
X4425 528 1 3994 539 4059 532 2 OAI22S $T=678900 376440 1 0 $X=678900 $Y=371020
X4426 3193 3269 3272 2 394 399 1 AO22 $T=549940 396600 0 0 $X=549940 $Y=396220
X4427 1294 1299 1262 1 2 1339 AO12 $T=239940 426840 0 0 $X=239940 $Y=426460
X4428 1320 1297 1316 1 2 1358 AO12 $T=243660 457080 1 0 $X=243660 $Y=451660
X4429 1370 1384 1396 1 2 1410 AO12 $T=257920 467160 1 0 $X=257920 $Y=461740
X4430 1322 1346 1414 1 2 59 AO12 $T=264120 396600 1 180 $X=260400 $Y=396220
X4431 1446 1453 1458 1 2 1465 AO12 $T=274660 487320 0 180 $X=270940 $Y=481900
X4432 1394 1289 1433 1 2 71 AO12 $T=271560 376440 1 0 $X=271560 $Y=371020
X4433 1485 1486 1481 1 2 1491 AO12 $T=282100 517560 0 180 $X=278380 $Y=512140
X4434 215 213 131 1 2 2033 AO12 $T=422220 366360 1 180 $X=418500 $Y=365980
X4435 2557 2584 258 1 2 2586 AO12 $T=453840 487320 1 0 $X=453840 $Y=481900
X4436 2971 3112 3125 1 2 3160 AO12 $T=528240 467160 1 0 $X=528240 $Y=461740
X4437 3186 340 3173 1 2 2841 AO12 $T=539400 376440 1 180 $X=535680 $Y=376060
X4438 3252 3182 3211 1 2 2798 AO12 $T=544360 386520 0 180 $X=540640 $Y=381100
X4439 3204 3208 3197 1 2 386 AO12 $T=544980 487320 1 180 $X=541260 $Y=486940
X4440 3238 3193 3201 1 2 3212 AO12 $T=545600 396600 1 180 $X=541880 $Y=396220
X4441 3158 3182 3212 1 2 3265 AO12 $T=543120 406680 1 0 $X=543120 $Y=401260
X4442 3225 3213 398 1 2 396 AO12 $T=553040 366360 1 180 $X=549320 $Y=365980
X4443 3734 3728 3719 1 2 3555 AO12 $T=625580 376440 1 180 $X=621860 $Y=376060
X4444 3873 3881 3876 1 2 3816 AO12 $T=652240 406680 1 180 $X=648520 $Y=406300
X4445 512 3920 3914 1 2 3711 AO12 $T=657820 386520 1 180 $X=654100 $Y=386140
X4446 3932 3984 3977 1 2 3940 AO12 $T=671460 436920 0 180 $X=667740 $Y=431500
X4447 1656 1644 2 1606 1 1662 AOI12HS $T=306280 386520 1 180 $X=301940 $Y=386140
X4448 1612 1651 2 1620 1 1655 AOI12HS $T=302560 376440 0 0 $X=302560 $Y=376060
X4449 1658 1646 2 1663 1 1696 AOI12HS $T=308140 436920 0 180 $X=303800 $Y=431500
X4450 1687 1683 2 1659 1 1665 AOI12HS $T=308140 497400 0 180 $X=303800 $Y=491980
X4451 1699 1677 2 1671 1 1654 AOI12HS $T=308760 457080 0 180 $X=304420 $Y=451660
X4452 1706 1677 2 1658 1 1739 AOI12HS $T=309380 436920 0 0 $X=309380 $Y=436540
X4453 1746 1731 2 1718 1 1690 AOI12HS $T=314960 487320 1 180 $X=310620 $Y=486940
X4454 1660 1709 2 1737 1 1755 AOI12HS $T=314340 396600 1 0 $X=314340 $Y=391180
X4455 1949 1906 2 1917 1 1965 AOI12HS $T=350920 507480 1 180 $X=346580 $Y=507100
X4456 1998 2019 2 1949 1 1912 AOI12HS $T=362080 507480 1 180 $X=357740 $Y=507100
X4457 2270 2235 2 2219 1 2014 AOI12HS $T=400520 507480 1 180 $X=396180 $Y=507100
X4458 2416 2418 2 2430 1 2453 AOI12HS $T=429040 507480 1 0 $X=429040 $Y=502060
X4459 2429 2446 2 2416 1 2449 AOI12HS $T=434000 497400 0 180 $X=429660 $Y=491980
X4460 2437 2476 2 2495 1 2510 AOI12HS $T=437100 426840 1 0 $X=437100 $Y=421420
X4461 2473 2477 2 2492 1 2468 AOI12HS $T=437100 507480 0 0 $X=437100 $Y=507100
X4462 2490 245 2 2514 1 2478 AOI12HS $T=438960 527640 0 0 $X=438960 $Y=527260
X4463 2627 2669 2 2661 1 2689 AOI12HS $T=466860 406680 1 0 $X=466860 $Y=401260
X4464 2724 2712 2 2750 1 2752 AOI12HS $T=478020 376440 0 0 $X=478020 $Y=376060
X4465 3131 2812 2 3092 1 3119 AOI12HS $T=531340 487320 0 180 $X=527000 $Y=481900
X4466 2816 3270 2 3311 1 3284 AOI12HS $T=554280 406680 0 0 $X=554280 $Y=406300
X4467 3476 3492 2 3507 1 3447 AOI12HS $T=587140 386520 1 0 $X=587140 $Y=381100
X4468 3521 3529 2 3539 1 3478 AOI12HS $T=592720 406680 0 0 $X=592720 $Y=406300
X4469 3525 3529 2 3540 1 3484 AOI12HS $T=592720 416760 1 0 $X=592720 $Y=411340
X4470 3509 3536 2 3530 1 3431 AOI12HS $T=593960 386520 0 0 $X=593960 $Y=386140
X4471 3522 3529 2 3547 1 3479 AOI12HS $T=593960 416760 0 0 $X=593960 $Y=416380
X4472 3528 3539 2 3576 1 3544 AOI12HS $T=598300 396600 0 0 $X=598300 $Y=396220
X4473 3547 3567 2 3595 1 3566 AOI12HS $T=601400 416760 0 0 $X=601400 $Y=416380
X4474 3569 3619 2 3631 1 3588 AOI12HS $T=606980 436920 1 0 $X=606980 $Y=431500
X4475 3619 3541 2 3650 1 3524 AOI12HS $T=609460 426840 0 0 $X=609460 $Y=426460
X4476 1207 2 1203 1261 1 AN2B1S $T=228160 436920 0 0 $X=228160 $Y=436540
X4477 1219 2 1231 1270 1 AN2B1S $T=229400 457080 1 0 $X=229400 $Y=451660
X4478 1268 2 1237 1284 1 AN2B1S $T=231260 396600 0 0 $X=231260 $Y=396220
X4479 1219 2 1241 1304 1 AN2B1S $T=236220 487320 1 0 $X=236220 $Y=481900
X4480 1319 2 1293 1362 1 AN2B1S $T=244900 507480 0 0 $X=244900 $Y=507100
X4481 51 2 1395 1427 1 AN2B1S $T=261020 527640 0 0 $X=261020 $Y=527260
X4482 67 2 68 1471 1 AN2B1S $T=269080 366360 0 0 $X=269080 $Y=365980
X4483 1459 2 68 1514 1 AN2B1S $T=277760 386520 0 0 $X=277760 $Y=386140
X4484 1476 2 1505 1510 1 AN2B1S $T=278380 416760 0 0 $X=278380 $Y=416380
X4485 1504 2 68 1519 1 AN2B1S $T=279620 406680 1 0 $X=279620 $Y=401260
X4486 51 2 1485 1525 1 AN2B1S $T=280240 527640 0 0 $X=280240 $Y=527260
X4487 1502 2 1505 1526 1 AN2B1S $T=280860 436920 0 0 $X=280860 $Y=436540
X4488 1520 2 1505 1533 1 AN2B1S $T=282100 426840 1 0 $X=282100 $Y=421420
X4489 1536 2 1505 1539 1 AN2B1S $T=284580 436920 0 0 $X=284580 $Y=436540
X4490 82 2 68 84 1 AN2B1S $T=287060 366360 0 0 $X=287060 $Y=365980
X4491 1550 2 1505 1577 1 AN2B1S $T=287680 436920 0 0 $X=287680 $Y=436540
X4492 1572 2 1578 1588 1 AN2B1S $T=292020 477240 1 0 $X=292020 $Y=471820
X4493 1583 2 1578 1575 1 AN2B1S $T=295740 467160 0 180 $X=292640 $Y=461740
X4494 1592 2 1578 1604 1 AN2B1S $T=295740 477240 1 0 $X=295740 $Y=471820
X4495 1717 2 1744 1769 1 AN2B1S $T=313100 517560 1 0 $X=313100 $Y=512140
X4496 1821 2 1744 1833 1 AN2B1S $T=326120 517560 1 0 $X=326120 $Y=512140
X4497 1858 2 1744 1924 1 AN2B1S $T=345340 517560 0 0 $X=345340 $Y=517180
X4498 1925 2 1744 1956 1 AN2B1S $T=349680 517560 0 0 $X=349680 $Y=517180
X4499 1927 2 1744 2093 1 AN2B1S $T=370140 517560 0 0 $X=370140 $Y=517180
X4500 2107 2 1744 2214 1 AN2B1S $T=384400 527640 1 0 $X=384400 $Y=522220
X4501 2161 2 184 2261 1 AN2B1S $T=394940 527640 0 0 $X=394940 $Y=527260
X4502 190 2 184 2279 1 AN2B1S $T=397420 537720 1 0 $X=397420 $Y=532300
X4503 2200 2 184 2297 1 AN2B1S $T=399900 527640 0 0 $X=399900 $Y=527260
X4504 228 2 2537 2464 1 AN2B1S $T=448260 426840 1 180 $X=445160 $Y=426460
X4505 2574 2 266 2598 1 AN2B1S $T=460660 406680 0 180 $X=457560 $Y=401260
X4506 284 2 273 2713 1 AN2B1S $T=471820 386520 0 0 $X=471820 $Y=386140
X4507 2812 2 2904 3048 1 AN2B1S $T=525140 497400 0 180 $X=522040 $Y=491980
X4508 1220 14 1 22 2 1256 OAI12HS $T=226300 537720 1 0 $X=226300 $Y=532300
X4509 1602 1591 1 1585 2 92 OAI12HS $T=298220 366360 1 180 $X=294500 $Y=365980
X4510 1607 1610 1 1598 2 1606 OAI12HS $T=300080 386520 1 180 $X=296360 $Y=386140
X4511 1640 1638 1 1657 2 1663 OAI12HS $T=301940 426840 0 0 $X=301940 $Y=426460
X4512 1666 1667 1 1645 2 1656 OAI12HS $T=306280 396600 1 180 $X=302560 $Y=396220
X4513 1649 1629 1 1641 2 1658 OAI12HS $T=306280 447000 0 180 $X=302560 $Y=441580
X4514 1679 1662 1 98 2 1661 OAI12HS $T=306900 386520 0 180 $X=303180 $Y=381100
X4515 1694 1690 1 1678 2 1659 OAI12HS $T=310000 487320 0 180 $X=306280 $Y=481900
X4516 1689 1702 1 1666 2 1722 OAI12HS $T=308140 406680 1 0 $X=308140 $Y=401260
X4517 1697 1702 1 1662 2 1651 OAI12HS $T=308760 386520 0 0 $X=308760 $Y=386140
X4518 1688 1702 1 1669 2 1709 OAI12HS $T=308760 396600 1 0 $X=308760 $Y=391180
X4519 1665 1711 1 1696 2 1710 OAI12HS $T=308760 436920 1 0 $X=308760 $Y=431500
X4520 1703 1716 1 1719 2 105 OAI12HS $T=312480 366360 0 0 $X=312480 $Y=365980
X4521 1623 1739 1 1640 2 1765 OAI12HS $T=313100 426840 0 0 $X=313100 $Y=426460
X4522 1715 1768 1 1690 2 1749 OAI12HS $T=318680 487320 1 180 $X=314960 $Y=486940
X4523 1797 1768 1 1778 2 1817 OAI12HS $T=322400 497400 0 0 $X=322400 $Y=497020
X4524 1721 1791 1 1871 2 128 OAI12HS $T=336040 376440 0 0 $X=336040 $Y=376060
X4525 1975 2014 1 1965 2 1687 OAI12HS $T=355260 507480 0 180 $X=351540 $Y=502060
X4526 2233 2202 1 2221 2 2219 OAI12HS $T=394940 507480 0 180 $X=391220 $Y=502060
X4527 2246 2256 1 2233 2 2224 OAI12HS $T=395560 507480 1 0 $X=395560 $Y=502060
X4528 2426 2438 1 2444 2 2437 OAI12HS $T=428420 426840 1 0 $X=428420 $Y=421420
X4529 2468 2456 1 2453 2 2270 OAI12HS $T=436480 507480 1 180 $X=432760 $Y=507100
X4530 2450 2478 1 2470 2 2477 OAI12HS $T=438960 527640 0 180 $X=435240 $Y=522220
X4531 2625 2592 1 2594 2 2603 OAI12HS $T=461280 457080 0 180 $X=457560 $Y=451660
X4532 2615 2510 1 2633 2 2627 OAI12HS $T=460040 416760 1 0 $X=460040 $Y=411340
X4533 2689 2693 1 2703 2 2712 OAI12HS $T=471820 406680 1 0 $X=471820 $Y=401260
X4534 2676 2706 1 2658 2 2709 OAI12HS $T=476780 447000 0 180 $X=473060 $Y=441580
X4535 2757 2752 1 2770 2 307 OAI12HS $T=482360 376440 0 0 $X=482360 $Y=376060
X4536 314 311 1 316 2 319 OAI12HS $T=489180 366360 0 0 $X=489180 $Y=365980
X4537 3254 3261 1 3203 2 3286 OAI12HS $T=555520 447000 0 180 $X=551800 $Y=441580
X4538 3364 3398 1 3325 2 3395 OAI12HS $T=574740 447000 0 180 $X=571020 $Y=441580
X4539 3445 434 1 3431 2 3438 OAI12HS $T=580940 386520 1 180 $X=577220 $Y=386140
X4540 3466 422 1 3447 2 3402 OAI12HS $T=584660 386520 0 180 $X=580940 $Y=381100
X4541 3500 434 1 3478 2 3483 OAI12HS $T=589620 406680 0 180 $X=585900 $Y=401260
X4542 3501 422 1 3479 2 3465 OAI12HS $T=589620 416760 1 180 $X=585900 $Y=416380
X4543 3512 422 1 3484 2 3472 OAI12HS $T=590860 416760 0 180 $X=587140 $Y=411340
X4544 3473 3470 1 3450 2 3513 OAI12HS $T=592720 447000 1 180 $X=589000 $Y=446620
X4545 3505 434 1 3524 2 3488 OAI12HS $T=590240 426840 1 0 $X=590240 $Y=421420
X4546 3511 422 1 3527 2 3487 OAI12HS $T=590860 396600 1 0 $X=590860 $Y=391180
X4547 3526 434 1 3537 2 3515 OAI12HS $T=592720 436920 1 0 $X=592720 $Y=431500
X4548 3558 3518 1 3458 2 3535 OAI12HS $T=597060 517560 0 180 $X=593340 $Y=512140
X4549 3519 3524 1 3544 2 3536 OAI12HS $T=593960 406680 1 0 $X=593960 $Y=401260
X4550 3563 3566 1 3580 2 3539 OAI12HS $T=599540 406680 0 0 $X=599540 $Y=406300
X4551 3579 422 1 3588 2 3599 OAI12HS $T=601400 426840 0 0 $X=601400 $Y=426460
X4552 3684 3673 1 3699 2 3690 OAI12HS $T=616900 447000 1 0 $X=616900 $Y=441580
X4553 3671 3606 1 3686 2 3650 OAI12HS $T=617520 426840 0 0 $X=617520 $Y=426460
X4554 479 486 1 480 2 3795 OAI12HS $T=637360 537720 0 180 $X=633640 $Y=532300
X4555 3790 3789 1 3817 2 3800 OAI12HS $T=637360 457080 0 0 $X=637360 $Y=456700
X4556 3839 3829 1 3766 2 3830 OAI12HS $T=643560 507480 1 180 $X=639840 $Y=507100
X4557 3741 3815 1 3852 2 3867 OAI12HS $T=649760 487320 0 180 $X=646040 $Y=481900
X4558 2880 2822 1 2892 2779 2910 2 MOAI1 $T=501580 426840 1 0 $X=501580 $Y=421420
X4559 3297 3316 1 3292 3190 3298 2 MOAI1 $T=559860 416760 1 180 $X=555520 $Y=416380
X4560 3337 3339 2992 1 2 OR2P $T=564200 416760 0 180 $X=560480 $Y=411340
X4561 2600 257 1 2 INV3 $T=461900 426840 0 0 $X=461900 $Y=426460
X4562 3104 3572 1 2 INV3 $T=599540 457080 0 0 $X=599540 $Y=456700
X4563 1560 2 1623 1579 1 1623 1646 1638 1202 ICV_22 $T=298840 436920 1 0 $X=298840 $Y=431500
X4564 1995 2 1983 2037 1 1995 2036 2045 1202 ICV_22 $T=362700 447000 1 0 $X=362700 $Y=441580
X4565 1969 2 2111 2098 1 2023 2117 2032 1202 ICV_22 $T=373240 477240 0 0 $X=373240 $Y=476860
X4566 2092 2 2085 2096 1 2106 2108 2128 1202 ICV_22 $T=373860 447000 0 0 $X=373860 $Y=446620
X4567 2091 2 2135 2096 1 2106 2141 2153 1202 ICV_22 $T=378200 447000 0 0 $X=378200 $Y=446620
X4568 2236 2 2234 186 1 2236 2254 2145 1202 ICV_22 $T=394320 406680 0 0 $X=394320 $Y=406300
X4569 185 2 2189 186 1 185 2252 182 1202 ICV_22 $T=394940 386520 1 0 $X=394940 $Y=381100
X4570 2245 2 2291 2061 1 2245 2263 1972 1202 ICV_22 $T=401760 467160 1 0 $X=401760 $Y=461740
X4571 2298 2 2300 2251 1 2298 2312 2288 1202 ICV_22 $T=404860 386520 1 0 $X=404860 $Y=381100
X4572 2637 2 2626 274 1 2659 2619 279 1202 ICV_22 $T=465000 527640 0 0 $X=465000 $Y=527260
X4573 2655 2 2678 2688 1 2665 2690 2658 1202 ICV_22 $T=469340 447000 1 0 $X=469340 $Y=441580
X4574 2519 2 2647 282 1 2547 2653 282 1202 ICV_22 $T=469960 467160 0 0 $X=469960 $Y=466780
X4575 288 2 2700 274 1 288 2708 271 1202 ICV_22 $T=471820 537720 1 0 $X=471820 $Y=532300
X4576 2778 2 2801 2814 1 2778 2818 2760 1202 ICV_22 $T=491040 497400 1 0 $X=491040 $Y=491980
X4577 3309 2 3308 3329 1 3338 3289 3349 1202 ICV_22 $T=559860 467160 1 0 $X=559860 $Y=461740
X4578 3317 2 3335 3305 1 3314 3347 3349 1202 ICV_22 $T=561100 477240 0 0 $X=561100 $Y=476860
X4579 3309 2 3553 3557 1 3305 3577 3408 1202 ICV_22 $T=597060 487320 1 0 $X=597060 $Y=481900
X4580 3418 2 3623 465 1 3617 3646 423 1202 ICV_22 $T=608220 517560 1 0 $X=608220 $Y=512140
X4581 3572 2 3676 3614 1 3614 3696 3636 1202 ICV_22 $T=615660 457080 0 0 $X=615660 $Y=456700
X4582 3103 231 2825 3104 1 2 QDFFRBP $T=528240 457080 0 0 $X=528240 $Y=456700
X4583 3235 231 3240 337 1 2 QDFFRBP $T=554900 537720 0 180 $X=542500 $Y=532300
X4584 3218 231 2825 3295 1 2 QDFFRBP $T=543740 467160 0 0 $X=543740 $Y=466780
X4585 3236 231 3288 365 1 2 QDFFRBP $T=545600 527640 1 0 $X=545600 $Y=522220
X4586 3245 231 3288 413 1 2 QDFFRBP $T=559240 527640 1 0 $X=559240 $Y=522220
X4587 5516 5680 1 2 BUF2CK $T=1021760 426840 0 0 $X=1021760 $Y=426460
X4588 3932 3941 3962 1 2 AN2T $T=658440 447000 1 0 $X=658440 $Y=441580
X4589 5100 1 5090 4661 2 810 ND3HT $T=901480 386520 1 180 $X=894040 $Y=386140
X4590 1246 1 1238 4 2 ND2P $T=228160 507480 1 180 $X=224440 $Y=507100
X4591 3299 1 3306 3249 2 ND2P $T=554900 386520 1 0 $X=554900 $Y=381100
X4592 247 2457 1 2523 2517 2544 2 MOAI1H $T=440200 467160 0 0 $X=440200 $Y=466780
X4593 1251 1260 1298 1 2 1312 HA1 $T=230020 406680 1 0 $X=230020 $Y=401260
X4594 1272 1279 37 1 2 1336 HA1 $T=234980 366360 0 0 $X=234980 $Y=365980
X4595 1274 1310 1364 1 2 1380 HA1 $T=243660 436920 0 0 $X=243660 $Y=436540
X4596 1311 1330 1388 1 2 1400 HA1 $T=248620 457080 1 0 $X=248620 $Y=451660
X4597 1281 1399 1430 1 2 1439 HA1 $T=257300 487320 0 0 $X=257300 $Y=486940
X4598 1391 1456 1487 1 2 1492 HA1 $T=269080 507480 0 0 $X=269080 $Y=507100
X4599 1464 1547 1580 1 2 1594 HA1 $T=287680 527640 0 0 $X=287680 $Y=527260
X4600 141 148 138 1 2 1926 HA1 $T=357120 537720 0 180 $X=349060 $Y=532300
X4601 154 2038 1948 1 2 1996 HA1 $T=365180 487320 1 180 $X=357120 $Y=486940
X4602 158 152 2044 1 2 2067 HA1 $T=358980 537720 1 0 $X=358980 $Y=532300
X4603 2057 2086 2043 1 2 2020 HA1 $T=372000 467160 1 180 $X=363940 $Y=466780
X4604 2085 2108 1966 1 2 2059 HA1 $T=375720 457080 0 180 $X=367660 $Y=451660
X4605 2127 2146 2110 1 2 2042 HA1 $T=381920 436920 0 180 $X=373860 $Y=431500
X4606 2117 2111 2133 1 2 2174 HA1 $T=376960 477240 0 0 $X=376960 $Y=476860
X4607 167 2188 2163 1 2 2138 HA1 $T=389980 467160 0 180 $X=381920 $Y=461740
X4608 173 2217 2177 1 2 2125 HA1 $T=391840 447000 1 180 $X=383780 $Y=446620
X4609 180 2193 2223 1 2 2226 HA1 $T=386880 426840 0 0 $X=386880 $Y=426460
X4610 181 2238 2151 1 2 2196 HA1 $T=396180 497400 0 180 $X=388120 $Y=491980
X4611 2277 2248 2228 1 2 2309 HA1 $T=399280 457080 1 0 $X=399280 $Y=451660
X4612 204 200 2318 1 2 2334 HA1 $T=401760 537720 1 0 $X=401760 $Y=532300
X4613 162 2293 2329 1 2 2357 HA1 $T=404240 457080 0 0 $X=404240 $Y=456700
X4614 2320 2255 2331 1 2 2342 HA1 $T=404860 487320 1 0 $X=404860 $Y=481900
X4615 192 2264 2338 1 2 2352 HA1 $T=404860 497400 0 0 $X=404860 $Y=497020
X4616 2253 2349 2367 1 2 2337 HA1 $T=423460 416760 1 180 $X=415400 $Y=416380
X4617 2341 2361 2167 1 2 2398 HA1 $T=416020 396600 0 0 $X=416020 $Y=396220
X4618 194 2242 2362 1 2 2370 HA1 $T=424700 447000 0 180 $X=416640 $Y=441580
X4619 2377 2383 2406 1 2 2403 HA1 $T=419740 487320 1 0 $X=419740 $Y=481900
X4620 2372 2427 2460 1 2 2440 HA1 $T=427800 426840 0 0 $X=427800 $Y=426460
X4621 2448 2419 237 1 2 2471 HA1 $T=428420 366360 0 0 $X=428420 $Y=365980
X4622 2479 2455 2486 1 2 2498 HA1 $T=432760 416760 1 0 $X=432760 $Y=411340
X4623 2497 2451 2513 1 2 2522 HA1 $T=435860 396600 1 0 $X=435860 $Y=391180
X4624 2585 2608 2575 1 2 2567 HA1 $T=459420 467160 0 180 $X=451360 $Y=461740
X4625 2647 2679 2638 1 2 2594 HA1 $T=469960 467160 1 180 $X=461900 $Y=466780
X4626 2717 2736 2701 1 2 2625 HA1 $T=480500 467160 0 180 $X=472440 $Y=461740
X4627 3274 3301 3259 1 2 2759 HA1 $T=556760 467160 0 180 $X=548700 $Y=461740
X4628 3154 3335 3302 1 2 3280 HA1 $T=562960 477240 0 180 $X=554900 $Y=471820
X4629 2982 3355 3383 1 2 3396 HA1 $T=564200 497400 1 0 $X=564200 $Y=491980
X4630 3371 3367 3391 1 2 3353 HA1 $T=566680 467160 1 0 $X=566680 $Y=461740
X4631 2941 3378 3407 1 2 3415 HA1 $T=568540 477240 0 0 $X=568540 $Y=476860
X4632 3543 3564 3531 1 2 3503 HA1 $T=600780 467160 0 180 $X=592720 $Y=461740
X4633 1205 6 1224 2 1 XOR2HS $T=220100 386520 0 0 $X=220100 $Y=386140
X4634 1206 6 1225 2 1 XOR2HS $T=220100 396600 0 0 $X=220100 $Y=396220
X4635 12 18 1212 2 1 XOR2HS $T=225680 426840 1 180 $X=220100 $Y=426460
X4636 7 9 1227 2 1 XOR2HS $T=220720 477240 1 0 $X=220720 $Y=471820
X4637 1217 13 1233 2 1 XOR2HS $T=221340 487320 0 0 $X=221340 $Y=486940
X4638 1230 18 1215 2 1 XOR2HS $T=227540 436920 1 180 $X=221960 $Y=436540
X4639 16 13 1239 2 1 XOR2HS $T=222580 487320 1 0 $X=222580 $Y=481900
X4640 1208 9 1259 2 1 XOR2HS $T=226920 477240 1 0 $X=226920 $Y=471820
X4641 25 29 1255 2 1 XOR2HS $T=233740 507480 1 180 $X=228160 $Y=507100
X4642 1305 29 1287 2 1 XOR2HS $T=239320 517560 0 180 $X=233740 $Y=512140
X4643 1305 52 1382 2 1 XOR2HS $T=250480 527640 1 0 $X=250480 $Y=522220
X4644 56 52 1383 2 1 XOR2HS $T=258540 527640 1 180 $X=252960 $Y=527260
X4645 1650 1655 1676 2 1 XOR2HS $T=303180 366360 0 0 $X=303180 $Y=365980
X4646 1611 1716 1742 2 1 XOR2HS $T=310620 376440 1 0 $X=310620 $Y=371020
X4647 1670 1654 1753 2 1 XOR2HS $T=311860 447000 1 0 $X=311860 $Y=441580
X4648 1621 1755 1771 2 1 XOR2HS $T=314340 386520 0 0 $X=314340 $Y=386140
X4649 1738 1702 1772 2 1 XOR2HS $T=314340 396600 0 0 $X=314340 $Y=396220
X4650 1781 1739 1804 2 1 XOR2HS $T=319920 426840 1 0 $X=319920 $Y=421420
X4651 1808 1768 1786 2 1 XOR2HS $T=325500 487320 1 180 $X=319920 $Y=486940
X4652 1913 1912 1890 2 1 XOR2HS $T=347200 497400 1 180 $X=341620 $Y=497020
X4653 2269 2256 2290 2 1 XOR2HS $T=399280 497400 0 0 $X=399280 $Y=497020
X4654 2428 2449 2472 2 1 XOR2HS $T=434620 497400 0 0 $X=434620 $Y=497020
X4655 2478 2504 2527 2 1 XOR2HS $T=440200 517560 0 0 $X=440200 $Y=517180
X4656 2563 2567 2542 2 1 XOR2HS $T=453220 457080 1 180 $X=447640 $Y=456700
X4657 2569 2571 2546 2 1 XOR2HS $T=454460 447000 0 180 $X=448880 $Y=441580
X4658 2572 261 2587 2 1 XOR2HS $T=451360 527640 0 0 $X=451360 $Y=527260
X4659 2624 2616 2600 2 1 XOR2HS $T=461900 426840 1 180 $X=456320 $Y=426460
X4660 2626 2619 2572 2 1 XOR2HS $T=461900 537720 0 180 $X=456320 $Y=532300
X4661 2587 265 2623 2 1 XOR2HS $T=456940 527640 0 0 $X=456940 $Y=527260
X4662 2616 2628 2607 2 1 XOR2HS $T=463760 436920 1 180 $X=458180 $Y=436540
X4663 2625 2592 2610 2 1 XOR2HS $T=463760 447000 1 180 $X=458180 $Y=446620
X4664 2580 2648 2634 2 1 XOR2HS $T=466860 517560 0 180 $X=461280 $Y=512140
X4665 2678 2674 2649 2 1 XOR2HS $T=469960 436920 1 180 $X=464380 $Y=436540
X4666 2665 2676 2655 2 1 XOR2HS $T=470580 447000 1 180 $X=465000 $Y=446620
X4667 287 283 2648 2 1 XOR2HS $T=471200 537720 0 180 $X=465620 $Y=532300
X4668 2668 2671 2686 2 1 XOR2HS $T=466860 507480 0 0 $X=466860 $Y=507100
X4669 2700 2696 2683 2 1 XOR2HS $T=474300 527640 1 180 $X=468720 $Y=527260
X4670 2676 2706 2688 2 1 XOR2HS $T=476160 447000 1 180 $X=470580 $Y=446620
X4671 2691 2683 2704 2 1 XOR2HS $T=470580 527640 1 0 $X=470580 $Y=522220
X4672 2699 2686 2719 2 1 XOR2HS $T=472440 507480 0 0 $X=472440 $Y=507100
X4673 2743 2708 2699 2 1 XOR2HS $T=481120 537720 0 180 $X=475540 $Y=532300
X4674 2715 2719 2741 2 1 XOR2HS $T=476160 517560 1 0 $X=476160 $Y=512140
X4675 2747 2674 2727 2 1 XOR2HS $T=482360 436920 1 180 $X=476780 $Y=436540
X4676 2738 2725 2756 2 1 XOR2HS $T=478640 527640 0 0 $X=478640 $Y=527260
X4677 2758 2761 2775 2 1 XOR2HS $T=481740 497400 0 0 $X=481740 $Y=497020
X4678 2733 2751 2780 2 1 XOR2HS $T=482360 517560 0 0 $X=482360 $Y=517180
X4679 2775 2776 2785 2 1 XOR2HS $T=484220 497400 1 0 $X=484220 $Y=491980
X4680 2777 2756 2787 2 1 XOR2HS $T=484840 527640 0 0 $X=484840 $Y=527260
X4681 2801 2794 2781 2 1 XOR2HS $T=491040 487320 0 180 $X=485460 $Y=481900
X4682 2787 2704 2804 2 1 XOR2HS $T=487320 527640 1 0 $X=487320 $Y=522220
X4683 2780 2791 2820 2 1 XOR2HS $T=490420 517560 0 0 $X=490420 $Y=517180
X4684 318 2819 2828 2 1 XOR2HS $T=491660 537720 1 0 $X=491660 $Y=532300
X4685 322 2828 2848 2 1 XOR2HS $T=493520 527640 0 0 $X=493520 $Y=527260
X4686 2832 2820 2850 2 1 XOR2HS $T=496620 517560 0 0 $X=496620 $Y=517180
X4687 2912 2915 2936 2 1 XOR2HS $T=505920 447000 0 0 $X=505920 $Y=446620
X4688 2936 3017 3064 2 1 XOR2HS $T=520800 457080 1 0 $X=520800 $Y=451660
X4689 3230 3229 2805 2 1 XOR2HS $T=546840 436920 0 180 $X=541260 $Y=431500
X4690 3220 3254 3234 2 1 XOR2HS $T=551180 447000 0 180 $X=545600 $Y=441580
X4691 3254 3261 3195 2 1 XOR2HS $T=551800 436920 1 180 $X=546220 $Y=436540
X4692 3279 3229 395 2 1 XOR2HS $T=553660 436920 0 180 $X=548080 $Y=431500
X4693 3328 3364 3374 2 1 XOR2HS $T=564820 447000 1 0 $X=564820 $Y=441580
X4694 3382 3379 414 2 1 XOR2HS $T=571020 426840 1 180 $X=565440 $Y=426460
X4695 3364 3398 3351 2 1 XOR2HS $T=575360 436920 1 180 $X=569780 $Y=436540
X4696 3382 3414 420 2 1 XOR2HS $T=577220 426840 1 180 $X=571640 $Y=426460
X4697 3452 434 3365 2 1 XOR2HS $T=583420 426840 0 180 $X=577840 $Y=421420
X4698 3453 3473 3485 2 1 XOR2HS $T=584040 447000 1 0 $X=584040 $Y=441580
X4699 3506 3502 445 2 1 XOR2HS $T=590860 436920 1 180 $X=585280 $Y=436540
X4700 3533 3506 452 2 1 XOR2HS $T=596440 436920 1 180 $X=590860 $Y=436540
X4701 3473 3470 3456 2 1 XOR2HS $T=597680 447000 0 180 $X=592100 $Y=441580
X4702 374 3542 3556 2 1 XOR2HS $T=594580 457080 1 0 $X=594580 $Y=451660
X4703 3558 3562 3586 2 1 XOR2HS $T=599540 517560 1 0 $X=599540 $Y=512140
X4704 3558 3518 3574 2 1 XOR2HS $T=600780 517560 0 0 $X=600780 $Y=517180
X4705 3601 3602 462 2 1 XOR2HS $T=604500 507480 1 0 $X=604500 $Y=502060
X4706 3684 3673 3718 2 1 XOR2HS $T=619380 436920 0 0 $X=619380 $Y=436540
X4707 3684 3716 3737 2 1 XOR2HS $T=621240 447000 0 0 $X=621240 $Y=446620
X4708 3651 3748 3757 2 1 XOR2HS $T=626200 436920 1 0 $X=626200 $Y=431500
X4709 479 3610 3788 2 1 XOR2HS $T=630540 527640 0 0 $X=630540 $Y=527260
X4710 3762 3780 487 2 1 XOR2HS $T=635500 447000 1 0 $X=635500 $Y=441580
X4711 479 486 3805 2 1 XOR2HS $T=637360 527640 0 0 $X=637360 $Y=527260
X4712 3790 3789 3828 2 1 XOR2HS $T=637980 457080 1 0 $X=637980 $Y=451660
X4713 3790 3835 3840 2 1 XOR2HS $T=641080 457080 0 0 $X=641080 $Y=456700
X4714 3762 3837 3849 2 1 XOR2HS $T=641700 447000 1 0 $X=641700 $Y=441580
X4715 3832 3794 3853 2 1 XOR2HS $T=642940 527640 0 0 $X=642940 $Y=527260
X4716 3839 3829 3871 2 1 XOR2HS $T=644800 497400 1 0 $X=644800 $Y=491980
X4717 3866 3843 500 2 1 XOR2HS $T=651620 467160 0 180 $X=646040 $Y=461740
X4718 3839 501 3883 2 1 XOR2HS $T=646660 507480 0 0 $X=646660 $Y=507100
X4719 3741 3815 3890 2 1 XOR2HS $T=647900 487320 0 0 $X=647900 $Y=486940
X4720 3866 3886 3897 2 1 XOR2HS $T=649140 477240 1 0 $X=649140 $Y=471820
X4721 504 499 3904 2 1 XOR2HS $T=650380 537720 1 0 $X=650380 $Y=532300
X4722 3741 3847 3912 2 1 XOR2HS $T=651620 487320 1 0 $X=651620 $Y=481900
X4723 3887 3906 3925 2 1 XOR2HS $T=652860 457080 1 0 $X=652860 $Y=451660
X4724 3900 3913 3941 2 1 XOR2HS $T=656580 517560 1 0 $X=656580 $Y=512140
X4725 504 515 3902 2 1 XOR2HS $T=656580 527640 0 0 $X=656580 $Y=527260
X4726 3655 3696 3717 1 2 3699 MAO222 $T=619380 457080 0 0 $X=619380 $Y=456700
X4727 3783 3749 3726 1 2 3815 MAO222 $T=634880 487320 0 0 $X=634880 $Y=486940
X4728 3781 3787 3747 1 2 3852 MAO222 $T=641080 487320 0 0 $X=641080 $Y=486940
X4729 10 1209 19 2 1 1242 XOR3 $T=239940 517560 1 180 $X=228780 $Y=517180
X4730 3655 3696 3717 2 1 3790 XOR3 $T=625580 457080 0 0 $X=625580 $Y=456700
X4731 3781 3787 3747 2 1 3839 XOR3 $T=633020 497400 1 0 $X=633020 $Y=491980
X4732 3783 3749 3726 2 1 3847 XOR3 $T=633640 487320 1 0 $X=633640 $Y=481900
X4733 2592 2653 2 2662 2638 1 2665 FA1 $T=455700 457080 0 0 $X=455700 $Y=456700
X4734 2658 2701 2 2710 2759 1 2676 FA1 $T=484840 457080 0 180 $X=469340 $Y=451660
X4735 2706 3280 2 3289 3216 1 3220 FA1 $T=542500 457080 1 0 $X=542500 $Y=451660
X4736 3203 3255 2 3350 3294 1 3254 FA1 $T=551800 447000 0 0 $X=551800 $Y=446620
X4737 3462 3403 2 3386 3409 1 3377 FA1 $T=584040 507480 0 180 $X=568540 $Y=502060
X4738 3325 3406 2 3381 3435 1 3364 FA1 $T=584660 447000 1 180 $X=569160 $Y=446620
X4739 3398 3474 2 3481 3439 1 3453 FA1 $T=575980 457080 1 0 $X=575980 $Y=451660
X4740 3458 3451 2 3534 3468 1 3558 FA1 $T=582800 517560 0 0 $X=582800 $Y=517180
X4741 3450 3489 2 3461 3552 1 3473 FA1 $T=583420 457080 0 0 $X=583420 $Y=456700
X4742 3470 3517 2 3462 3482 1 3562 FA1 $T=584660 507480 1 0 $X=584660 $Y=502060
X4743 3518 3433 2 458 454 1 3610 FA1 $T=591480 527640 0 0 $X=591480 $Y=527260
X4744 3640 3623 2 405 3624 1 3746 FA1 $T=610700 517560 0 0 $X=610700 $Y=517180
X4745 3741 3770 2 3638 3725 1 3817 FA1 $T=625580 477240 0 0 $X=625580 $Y=476860
X4746 3766 3785 2 3727 3740 1 3829 FA1 $T=631160 517560 1 0 $X=631160 $Y=512140
X4747 3770 3733 2 3126 3769 1 3865 FA1 $T=631780 477240 1 0 $X=631780 $Y=471820
X4748 3835 3786 2 3724 3865 1 3789 FA1 $T=651000 467160 1 180 $X=635500 $Y=466780
X4749 546 4025 2 4008 4066 1 3731 FA1 $T=686960 396600 0 180 $X=671460 $Y=391180
X4750 4026 3937 2 3860 4007 1 4076 FA1 $T=676420 406680 1 0 $X=676420 $Y=401260
X4751 561 4061 2 4092 4093 1 4066 FA1 $T=699980 376440 1 180 $X=684480 $Y=376060
X4752 3340 399 2 1 3187 3334 410 3365 3361 3346 3360 1202 ICV_24 $T=565440 376440 1 180 $X=561100 $Y=376060
X4753 4376 4356 2 1 4360 4359 4159 4152 4383 621 4374 1202 ICV_24 $T=748340 396600 1 180 $X=744000 $Y=396220
X4754 4439 4430 2 1 4434 4407 4410 4412 4457 4422 4471 1202 ICV_24 $T=766320 416760 0 180 $X=761980 $Y=411340
X4755 3907 4524 2 1 4504 4399 4316 4530 4512 3784 3857 1202 ICV_24 $T=776860 487320 0 180 $X=772520 $Y=481900
X4756 4509 4513 2 1 4517 4459 651 4306 4525 4479 4419 1202 ICV_24 $T=778720 507480 0 180 $X=774380 $Y=502060
X4757 3621 654 2 1 4531 4496 653 655 4521 3551 3587 1202 ICV_24 $T=782440 527640 1 180 $X=778100 $Y=527260
X4758 773 775 2 1 4934 722 776 779 4857 780 782 1202 ICV_24 $T=868620 537720 0 180 $X=864280 $Y=532300
X4759 5203 783 2 1 831 833 5153 4891 5202 838 843 1202 ICV_24 $T=919460 376440 0 180 $X=915120 $Y=371020
X4760 5290 5048 2 1 5281 5207 873 871 5193 5314 5270 1202 ICV_24 $T=938680 497400 0 180 $X=934340 $Y=491980
X4761 5722 5571 2 1 5695 5668 5573 5613 5726 5740 5717 1202 ICV_24 $T=1032300 406680 1 180 $X=1027960 $Y=406300
X4762 5776 5466 2 1 5755 5765 5709 5787 5784 1060 5772 1202 ICV_24 $T=1045320 447000 1 180 $X=1040980 $Y=446620
X4763 5832 5810 2 1 5814 1065 5760 5680 5830 5826 5818 1202 ICV_24 $T=1055860 426840 0 180 $X=1051520 $Y=421420
X4764 1073 5681 2 1 5815 5765 1047 5787 5823 5835 5844 1202 ICV_24 $T=1055860 447000 1 180 $X=1051520 $Y=446620
X4765 5843 5836 2 1 5840 5859 1007 5641 5877 5885 5820 1202 ICV_24 $T=1065160 517560 1 180 $X=1060820 $Y=517180
X4766 5994 5858 2 1 5947 5911 5749 5829 5982 5958 6009 1202 ICV_24 $T=1090580 497400 0 180 $X=1086240 $Y=491980
X4767 5975 5854 2 1 5977 5969 5760 5680 5970 6008 5955 1202 ICV_24 $T=1091200 416760 1 180 $X=1086860 $Y=416380
X4768 4161 2 1 4410 BUF3 $T=749580 416760 1 0 $X=749580 $Y=411340
X4769 880 2 1 871 BUF3 $T=944260 537720 0 180 $X=940540 $Y=532300
X4770 1941 1952 1959 1 2 150 AN3S $T=350300 376440 1 0 $X=350300 $Y=371020
X4771 4409 4707 4710 1 2 694 AN3S $T=815920 436920 1 0 $X=815920 $Y=431500
X4772 4285 4783 4791 1 2 719 AN3S $T=835140 487320 0 0 $X=835140 $Y=486940
X4773 3572 1 465 2 BUF4CK $T=611940 507480 1 0 $X=611940 $Y=502060
X4774 2400 2475 239 2025 2 2485 1 AOI13HS $T=435860 406680 1 0 $X=435860 $Y=401260
X4775 2730 2803 2788 2789 2 258 1 AOI13HS $T=492900 436920 0 180 $X=489180 $Y=431500
X4776 3224 3267 3117 3122 2 3282 1 AOI13HS $T=549940 507480 1 0 $X=549940 $Y=502060
X4777 450 430 1 2 BUF6 $T=589620 487320 1 0 $X=589620 $Y=481900
X4778 3920 521 1 2 BUF6 $T=659680 386520 1 0 $X=659680 $Y=381100
X4779 4407 637 1 2 BUF6 $T=756400 386520 0 0 $X=756400 $Y=386140
X4780 637 784 1 2 BUF6 $T=872340 366360 0 0 $X=872340 $Y=365980
X4781 107 1801 1596 1823 2 1 MXL2HS $T=323020 457080 1 0 $X=323020 $Y=451660
X4782 117 1801 1614 1818 2 1 MXL2HS $T=323640 436920 0 0 $X=323640 $Y=436540
X4783 108 1801 1673 1831 2 1 MXL2HS $T=324260 467160 1 0 $X=324260 $Y=461740
X4784 1796 1578 1794 1847 2 1 MXL2HS $T=326740 477240 0 0 $X=326740 $Y=476860
X4785 1721 122 1576 1839 2 1 MXL2HS $T=334800 376440 1 180 $X=329220 $Y=376060
X4786 1840 1801 1622 1857 2 1 MXL2HS $T=329220 426840 0 0 $X=329220 $Y=426460
X4787 1844 122 124 1867 2 1 MXL2HS $T=332320 366360 0 0 $X=332320 $Y=365980
X4788 125 1837 1736 1854 2 1 MXL2HS $T=337900 477240 1 180 $X=332320 $Y=476860
X4789 1828 1860 1571 1872 2 1 MXL2HS $T=334180 386520 0 0 $X=334180 $Y=386140
X4790 1803 1860 1595 1877 2 1 MXL2HS $T=334800 416760 0 0 $X=334800 $Y=416380
X4791 1845 1860 1681 1878 2 1 MXL2HS $T=335420 416760 1 0 $X=335420 $Y=411340
X4792 1791 1860 1587 1907 2 1 MXL2HS $T=340380 396600 0 0 $X=340380 $Y=396220
X4793 1815 1860 1619 1908 2 1 MXL2HS $T=340380 406680 0 0 $X=340380 $Y=406300
X4794 1862 1837 1940 1955 2 1 MXL2HS $T=347200 497400 0 0 $X=347200 $Y=497020
X4795 2212 1837 2008 2144 2 1 MXL2HS $T=391220 497400 1 180 $X=385640 $Y=497020
X4796 2299 2280 2131 2243 2 1 MXL2HS $T=406100 477240 0 180 $X=400520 $Y=471820
X4797 2372 212 2358 2318 2 1 MXL2HS $T=418500 527640 1 180 $X=412920 $Y=527260
X4798 2374 2280 2346 2323 2 1 MXL2HS $T=419740 497400 0 180 $X=414160 $Y=491980
X4799 2375 2347 2360 2352 2 1 MXL2HS $T=419740 507480 0 180 $X=414160 $Y=502060
X4800 2380 2347 2368 2363 2 1 MXL2HS $T=420360 507480 1 180 $X=414780 $Y=507100
X4801 2399 2280 2295 2353 2 1 MXL2HS $T=424080 477240 0 180 $X=418500 $Y=471820
X4802 2402 2280 2178 2379 2 1 MXL2HS $T=424700 467160 0 180 $X=419120 $Y=461740
X4803 2411 2280 2332 2389 2 1 MXL2HS $T=426560 497400 0 180 $X=420980 $Y=491980
X4804 1 2 1132 ANTENNA $T=1125920 386520 1 0 $X=1125920 $Y=381100
X4805 477 1 2 484 3707 3736 3742 3759 1202 ICV_30 $T=620000 527640 1 0 $X=620000 $Y=522220
X4806 3947 1 2 3996 3927 3955 3961 3966 1202 ICV_30 $T=657200 497400 1 0 $X=657200 $Y=491980
X4807 631 1 2 638 4373 4396 623 630 1202 ICV_30 $T=747100 366360 0 0 $X=747100 $Y=365980
X4808 4499 1 2 4510 4490 4537 4527 4554 1202 ICV_30 $T=779340 386520 1 0 $X=779340 $Y=381100
X4809 4750 1 2 4749 4612 4655 4690 4697 1202 ICV_30 $T=819640 416760 1 0 $X=819640 $Y=411340
X4810 4929 1 2 4968 4836 4920 4905 4944 1202 ICV_30 $T=861800 457080 1 0 $X=861800 $Y=451660
X4811 5177 1 2 5178 5078 5105 5080 5134 1202 ICV_30 $T=903340 477240 0 0 $X=903340 $Y=476860
X4812 838 1 2 5203 793 5053 5142 5180 1202 ICV_30 $T=908920 366360 0 0 $X=908920 $Y=365980
X4813 993 1 2 999 5532 5529 985 992 1202 ICV_30 $T=992000 527640 1 0 $X=992000 $Y=522220
X4814 5633 1 2 5631 995 1002 5606 5621 1202 ICV_30 $T=1002540 376440 0 0 $X=1002540 $Y=376060
X4815 5868 1 2 5867 5793 5811 5846 5864 1202 ICV_30 $T=1053380 507480 1 0 $X=1053380 $Y=502060
X4816 5941 1 2 5906 5860 5888 5828 5839 1202 ICV_30 $T=1071980 386520 0 0 $X=1071980 $Y=386140
X4817 6030 1 2 6048 6021 6015 6020 6034 1202 ICV_30 $T=1095540 467160 0 0 $X=1095540 $Y=466780
X4818 6064 1 2 6086 6018 6022 6009 5994 1202 ICV_30 $T=1095540 507480 1 0 $X=1095540 $Y=502060
X4819 1128 1 2 1133 6105 6106 6088 6120 1202 ICV_30 $T=1112280 436920 1 0 $X=1112280 $Y=431500
X4820 6045 1 2 6072 6108 6111 5874 5929 1202 ICV_30 $T=1112900 406680 1 0 $X=1112900 $Y=401260
X4821 1130 1 2 1136 1120 6113 1127 1129 1202 ICV_30 $T=1114760 366360 0 0 $X=1114760 $Y=365980
X4822 1131 1 2 1137 6085 6097 6016 6040 1202 ICV_30 $T=1114760 497400 1 0 $X=1114760 $Y=491980
X4823 4195 4154 4184 568 4134 1 2 AN4B1 $T=709280 426840 0 180 $X=703700 $Y=421420
X4824 4251 4264 4282 588 4284 1 2 AN4B1 $T=726020 406680 1 0 $X=726020 $Y=401260
X4825 5501 5490 5399 4141 5483 1 2 AN4B1 $T=987040 467160 0 180 $X=981460 $Y=461740
X4826 5499 5508 5221 4282 5518 1 2 AN4B1 $T=986420 406680 1 0 $X=986420 $Y=401260
X4827 557 1 2 4242 BUF8CK $T=715480 467160 0 0 $X=715480 $Y=466780
X4828 2537 2546 1 2554 2 AN2S $T=446400 447000 1 0 $X=446400 $Y=441580
X4829 2649 273 1 2672 2 AN2S $T=465620 426840 1 0 $X=465620 $Y=421420
X4830 301 2805 1 2786 2 AN2S $T=490420 376440 1 0 $X=490420 $Y=371020
X4831 492 3853 1 3863 2 AN2S $T=645420 376440 1 0 $X=645420 $Y=371020
X4832 3916 3925 1 3942 2 AN2S $T=657820 447000 0 0 $X=657820 $Y=446620
X4833 3909 3932 1 2 INV4 $T=656580 517560 0 0 $X=656580 $Y=517180
X4834 3771 3694 1 3694 494 3778 2 MOAI1HP $T=632400 507480 1 0 $X=632400 $Y=502060
X4835 3278 3276 1 3270 3108 2816 2 OAI22H $T=554900 416760 0 180 $X=547460 $Y=411340
X4836 3298 3356 1 3327 3376 3324 2 OAI22H $T=563580 406680 0 0 $X=563580 $Y=406300
X4837 3319 408 3307 1 2 XNR2H $T=556760 426840 0 0 $X=556760 $Y=426460
X4838 3049 3042 3081 2 3098 1 3142 AO112 $T=527620 497400 1 0 $X=527620 $Y=491980
X4839 3235 3204 2999 2 3251 1 3262 AO112 $T=545600 487320 0 0 $X=545600 $Y=486940
X4840 2946 3135 3076 3122 3107 372 1 2 3090 AO222 $T=533200 517560 1 180 $X=527000 $Y=517180
X4841 2971 3069 3113 374 3134 3041 1 2 3103 AO222 $T=527620 477240 1 0 $X=527620 $Y=471820
X4842 2847 3091 3041 3113 3134 3020 1 2 3164 AO222 $T=529480 477240 0 0 $X=529480 $Y=476860
X4843 2847 3055 3020 3113 3134 3177 1 2 3199 AO222 $T=533820 477240 1 0 $X=533820 $Y=471820
X4844 3105 3135 3166 3122 3107 3185 1 2 3192 AO222 $T=534440 517560 0 0 $X=534440 $Y=517180
X4845 3070 3135 3214 3122 3107 3228 1 2 3236 AO222 $T=540640 517560 0 0 $X=540640 $Y=517180
X4846 2990 3135 3219 3122 3107 3095 1 2 3245 AO222 $T=541260 517560 1 0 $X=541260 $Y=512140
X4847 3078 2802 2918 359 355 2938 2 1 2907 OA222S $T=524520 406680 0 180 $X=518940 $Y=401260
X4848 2779 231 2783 2 1 2792 QDFFRBS $T=484840 416760 0 0 $X=484840 $Y=416380
X4849 1701 1710 2 106 1661 1 AOI12H $T=310000 386520 1 0 $X=310000 $Y=381100
.ENDS
***************************************
.SUBCKT AN3B2S I1 B2 VCC B1 GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR3 I3 I2 I1 VCC GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV2CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MOAI1HT B1 B2 GND A1 O A2 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2B1 B1 I1 GND VCC O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI222S C1 C2 GND B1 B2 VCC A1 O A2
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2T I2 I1 GND O VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI12HP B2 B1 VCC O A1 GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI12H B2 B1 GND A1 O VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI12HP B2 B1 GND A1 O VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR2T O I2 GND I1 VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI12HT B2 B1 GND A1 O VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540
+ 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560
+ 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580
+ 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640
+ 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660
+ 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680
+ 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700
+ 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720
+ 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740
+ 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760
+ 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780
+ 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800
+ 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820
+ 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840
+ 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860
+ 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880
+ 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900
+ 901 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920
+ 921 922 923 924 925 926 927 928 929 930 931 932 933 934 935 936 937 938 939 940
+ 941 942 943 944 945 946 947 948 949 950 951 952 953 954 955 956 957 958 959 960
+ 961 962 963 964 965 966 967 968 969 970 971 972 973 974 975 976 977 978 979 980
+ 981 982 983 984 985 986 987 988 989 990 991 992 993 994 995 996 997 998 999 1000
+ 1001 1002 1003 1004 1005 1006 1007 1008 1009 1010 1011 1012 1013 1014 1015 1016 1017 1018 1019 1020
+ 1021 1022 1023 1024 1025 1026 1027 1028 1029 1030 1031 1032 1033 1034 1035 1036 1037 1038 1039 1040
+ 1041 1042 1043 1044 1045 1046 1047 1048 1049 1050 1051 1052 1053 1054 1055 1056 1057 1058 1070
** N=3804 EP=1059 IP=18566 FDC=0
X0 1057 3803 3803 3803 2954 3803 1058 YA2GSD $T=1349740 304020 0 90 $X=1210240 $Y=306870
X1 1073 2 3 1 INV1S $T=221340 265560 1 180 $X=220100 $Y=265180
X2 1071 2 6 1 INV1S $T=220100 295800 1 0 $X=220100 $Y=290380
X3 1072 2 1083 1 INV1S $T=221960 315960 0 0 $X=221960 $Y=315580
X4 1075 2 1082 1 INV1S $T=221960 346200 0 0 $X=221960 $Y=345820
X5 1094 2 1087 1 INV1S $T=225680 285720 0 180 $X=224440 $Y=280300
X6 1090 2 1101 1 INV1S $T=226920 356280 0 0 $X=226920 $Y=355900
X7 1071 2 1091 1 INV1S $T=228780 305880 0 180 $X=227540 $Y=300460
X8 1107 2 1108 1 INV1S $T=231260 305880 0 180 $X=230020 $Y=300460
X9 16 2 1071 1 INV1S $T=230020 305880 0 0 $X=230020 $Y=305500
X10 1105 2 1109 1 INV1S $T=230640 336120 1 0 $X=230640 $Y=330700
X11 1103 2 1116 1 INV1S $T=231880 275640 0 0 $X=231880 $Y=275260
X12 1083 2 1117 1 INV1S $T=233120 305880 0 0 $X=233120 $Y=305500
X13 21 2 26 1 INV1S $T=238700 265560 0 180 $X=237460 $Y=260140
X14 21 2 1142 1 INV1S $T=239940 265560 0 0 $X=239940 $Y=265180
X15 1142 2 1114 1 INV1S $T=241800 275640 1 180 $X=240560 $Y=275260
X16 1130 2 1145 1 INV1S $T=241800 305880 0 0 $X=241800 $Y=305500
X17 1142 2 34 1 INV1S $T=242420 265560 0 0 $X=242420 $Y=265180
X18 1083 2 1140 1 INV1S $T=245520 315960 1 180 $X=244280 $Y=315580
X19 1083 2 1155 1 INV1S $T=245520 315960 1 0 $X=245520 $Y=310540
X20 1163 2 1158 1 INV1S $T=248000 275640 0 180 $X=246760 $Y=270220
X21 1155 2 1166 1 INV1S $T=246760 315960 1 0 $X=246760 $Y=310540
X22 1149 2 1157 1 INV1S $T=246760 346200 1 0 $X=246760 $Y=340780
X23 1120 2 1163 1 INV1S $T=247380 265560 0 0 $X=247380 $Y=265180
X24 1163 2 43 1 INV1S $T=248620 265560 0 0 $X=248620 $Y=265180
X25 1137 2 58 1 INV1S $T=258540 275640 0 0 $X=258540 $Y=275260
X26 1134 2 61 1 INV1S $T=259780 265560 1 0 $X=259780 $Y=260140
X27 63 2 57 1 INV1S $T=266600 265560 0 180 $X=265360 $Y=260140
X28 1154 2 1221 1 INV1S $T=265360 265560 0 0 $X=265360 $Y=265180
X29 1136 2 64 1 INV1S $T=265360 275640 1 0 $X=265360 $Y=270220
X30 1209 2 1216 1 INV1S $T=266600 295800 0 0 $X=266600 $Y=295420
X31 1235 2 1223 1 INV1S $T=268460 265560 0 180 $X=267220 $Y=260140
X32 1196 2 1229 1 INV1S $T=267220 305880 1 0 $X=267220 $Y=300460
X33 1333 2 1306 1 INV1S $T=306900 326040 1 180 $X=305660 $Y=325660
X34 1333 2 92 1 INV1S $T=309380 315960 0 180 $X=308140 $Y=310540
X35 1322 2 1335 1 INV1S $T=309380 366360 0 180 $X=308140 $Y=360940
X36 1346 2 1350 1 INV1S $T=309380 336120 0 0 $X=309380 $Y=335740
X37 1352 2 1377 1 INV1S $T=314960 346200 0 0 $X=314960 $Y=345820
X38 1401 2 1394 1 INV1S $T=323020 326040 1 180 $X=321780 $Y=325660
X39 1412 2 1419 1 INV1S $T=324880 315960 0 0 $X=324880 $Y=315580
X40 1415 2 1422 1 INV1S $T=325500 295800 1 0 $X=325500 $Y=290380
X41 1405 2 1418 1 INV1S $T=326740 305880 0 180 $X=325500 $Y=300460
X42 1421 2 1424 1 INV1S $T=326120 285720 0 0 $X=326120 $Y=285340
X43 1429 2 1433 1 INV1S $T=330460 265560 0 180 $X=329220 $Y=260140
X44 1417 2 1440 1 INV1S $T=329840 275640 1 0 $X=329840 $Y=270220
X45 104 2 1333 1 INV1S $T=331080 336120 0 180 $X=329840 $Y=330700
X46 1333 2 1457 1 INV1S $T=333560 315960 1 0 $X=333560 $Y=310540
X47 1409 2 1470 1 INV1S $T=339140 346200 1 180 $X=337900 $Y=345820
X48 1478 2 1482 1 INV1S $T=340380 356280 0 0 $X=340380 $Y=355900
X49 1487 2 1480 1 INV1S $T=342240 295800 1 180 $X=341000 $Y=295420
X50 1464 2 1485 1 INV1S $T=341000 336120 0 0 $X=341000 $Y=335740
X51 1462 2 1486 1 INV1S $T=342860 356280 0 180 $X=341620 $Y=350860
X52 114 2 116 1 INV1S $T=345960 366360 1 0 $X=345960 $Y=360940
X53 1448 2 1516 1 INV1S $T=350300 346200 1 0 $X=350300 $Y=340780
X54 112 2 1517 1 INV1S $T=351540 336120 1 0 $X=351540 $Y=330700
X55 119 2 115 1 INV1S $T=352160 356280 1 0 $X=352160 $Y=350860
X56 121 2 1521 1 INV1S $T=352780 326040 0 0 $X=352780 $Y=325660
X57 128 2 1519 1 INV1S $T=354020 336120 1 180 $X=352780 $Y=335740
X58 125 2 1520 1 INV1S $T=354640 326040 0 180 $X=353400 $Y=320620
X59 129 2 1526 1 INV1S $T=354020 366360 1 0 $X=354020 $Y=360940
X60 136 2 1536 1 INV1S $T=358980 366360 1 0 $X=358980 $Y=360940
X61 123 2 139 1 INV1S $T=360220 366360 1 0 $X=360220 $Y=360940
X62 1527 2 1552 1 INV1S $T=368280 305880 0 180 $X=367040 $Y=300460
X63 1512 2 1607 1 INV1S $T=382540 295800 1 0 $X=382540 $Y=290380
X64 1647 2 165 1 INV1S $T=391220 305880 0 0 $X=391220 $Y=305500
X65 1527 2 1652 1 INV1S $T=391840 295800 0 0 $X=391840 $Y=295420
X66 1647 2 1660 1 INV1S $T=397420 295800 0 180 $X=396180 $Y=290380
X67 1628 2 171 1 INV1S $T=396800 356280 0 0 $X=396800 $Y=355900
X68 161 2 1647 1 INV1S $T=400520 285720 0 180 $X=399280 $Y=280300
X69 173 2 177 1 INV1S $T=399280 366360 1 0 $X=399280 $Y=360940
X70 173 2 1668 1 INV1S $T=400520 326040 1 0 $X=400520 $Y=320620
X71 173 2 1677 1 INV1S $T=402380 356280 1 0 $X=402380 $Y=350860
X72 1694 2 1659 1 INV1S $T=404240 326040 1 180 $X=403000 $Y=325660
X73 182 2 1619 1 INV1S $T=405480 275640 1 180 $X=404240 $Y=275260
X74 1694 2 183 1 INV1S $T=406100 326040 0 0 $X=406100 $Y=325660
X75 170 2 1694 1 INV1S $T=407960 295800 0 180 $X=406720 $Y=290380
X76 1697 2 1713 1 INV1S $T=413540 265560 1 0 $X=413540 $Y=260140
X77 144 2 209 1 INV1S $T=425940 356280 1 0 $X=425940 $Y=350860
X78 208 2 145 1 INV1S $T=429040 356280 1 0 $X=429040 $Y=350860
X79 211 2 192 1 INV1S $T=429040 356280 0 0 $X=429040 $Y=355900
X80 1745 2 1748 1 INV1S $T=429660 315960 1 0 $X=429660 $Y=310540
X81 218 2 201 1 INV1S $T=434620 366360 0 180 $X=433380 $Y=360940
X82 218 2 1779 1 INV1S $T=436480 346200 1 0 $X=436480 $Y=340780
X83 198 2 220 1 INV1S $T=437720 366360 0 180 $X=436480 $Y=360940
X84 1863 2 1854 1 INV1S $T=467480 336120 1 180 $X=466240 $Y=335740
X85 243 2 1863 1 INV1S $T=468100 336120 0 0 $X=468100 $Y=335740
X86 1863 2 1883 1 INV1S $T=474300 346200 0 0 $X=474300 $Y=345820
X87 258 2 1889 1 INV1S $T=477400 285720 1 180 $X=476160 $Y=285340
X88 259 2 1868 1 INV1S $T=477400 346200 0 180 $X=476160 $Y=340780
X89 266 2 1886 1 INV1S $T=481120 346200 0 180 $X=479880 $Y=340780
X90 269 2 1914 1 INV1S $T=482980 366360 1 0 $X=482980 $Y=360940
X91 258 2 1890 1 INV1S $T=484840 326040 1 180 $X=483600 $Y=325660
X92 265 2 1902 1 INV1S $T=485460 336120 0 180 $X=484220 $Y=330700
X93 271 2 1936 1 INV1S $T=490420 366360 1 0 $X=490420 $Y=360940
X94 1956 2 1959 1 INV1S $T=498480 346200 1 0 $X=498480 $Y=340780
X95 1969 2 1972 1 INV1S $T=504680 336120 1 180 $X=503440 $Y=335740
X96 1970 2 1978 1 INV1S $T=504060 346200 0 0 $X=504060 $Y=345820
X97 1974 2 1996 1 INV1S $T=509640 336120 1 0 $X=509640 $Y=330700
X98 1981 2 2024 1 INV1S $T=514600 336120 0 0 $X=514600 $Y=335740
X99 2018 2 2029 1 INV1S $T=516460 336120 1 0 $X=516460 $Y=330700
X100 2041 2 2060 1 INV1S $T=523280 326040 1 0 $X=523280 $Y=320620
X101 2073 2 2088 1 INV1S $T=530100 326040 1 0 $X=530100 $Y=320620
X102 312 2 2091 1 INV1S $T=533200 356280 0 0 $X=533200 $Y=355900
X103 314 2 2092 1 INV1S $T=535680 356280 1 180 $X=534440 $Y=355900
X104 2097 2 2107 1 INV1S $T=536300 326040 1 0 $X=536300 $Y=320620
X105 2103 2 2106 1 INV1S $T=537540 315960 0 0 $X=537540 $Y=315580
X106 2094 2 2120 1 INV1S $T=538160 315960 1 0 $X=538160 $Y=310540
X107 322 2 2114 1 INV1S $T=541260 356280 0 180 $X=540020 $Y=350860
X108 2143 2 2148 1 INV1S $T=546220 305880 0 0 $X=546220 $Y=305500
X109 2131 2 2154 1 INV1S $T=546840 326040 1 0 $X=546840 $Y=320620
X110 2136 2 2153 1 INV1S $T=547460 305880 1 0 $X=547460 $Y=300460
X111 2161 2 2151 1 INV1S $T=549940 295800 1 180 $X=548700 $Y=295420
X112 333 2 2163 1 INV1S $T=548700 305880 1 0 $X=548700 $Y=300460
X113 2157 2 2141 1 INV1S $T=549320 315960 0 0 $X=549320 $Y=315580
X114 2198 2 2161 1 INV1S $T=559860 275640 1 180 $X=558620 $Y=275260
X115 346 2 2195 1 INV1S $T=558620 366360 1 0 $X=558620 $Y=360940
X116 2198 2 2187 1 INV1S $T=559860 275640 0 0 $X=559860 $Y=275260
X117 1987 2 2230 1 INV1S $T=564200 285720 1 0 $X=564200 $Y=280300
X118 357 2 2213 1 INV1S $T=566680 295800 0 180 $X=565440 $Y=290380
X119 2230 2 361 1 INV1S $T=566680 285720 1 0 $X=566680 $Y=280300
X120 2228 2 2229 1 INV1S $T=567920 295800 0 180 $X=566680 $Y=290380
X121 2230 2 2239 1 INV1S $T=567920 285720 1 0 $X=567920 $Y=280300
X122 2233 2 2209 1 INV1S $T=569160 295800 0 180 $X=567920 $Y=290380
X123 2040 2 1772 1 INV1S $T=571640 346200 0 0 $X=571640 $Y=345820
X124 2240 2 2264 1 INV1S $T=577220 305880 1 0 $X=577220 $Y=300460
X125 2257 2 2266 1 INV1S $T=577840 275640 0 0 $X=577840 $Y=275260
X126 259 2 2272 1 INV1S $T=578460 346200 1 0 $X=578460 $Y=340780
X127 2250 2 2279 1 INV1S $T=580940 295800 0 0 $X=580940 $Y=295420
X128 2275 2 2269 1 INV1S $T=582800 326040 1 180 $X=581560 $Y=325660
X129 2272 2 384 1 INV1S $T=581560 346200 1 0 $X=581560 $Y=340780
X130 379 2 2292 1 INV1S $T=587760 295800 0 0 $X=587760 $Y=295420
X131 2311 2 2308 1 INV1S $T=592100 315960 1 180 $X=590860 $Y=315580
X132 2301 2 2306 1 INV1S $T=593340 285720 1 180 $X=592100 $Y=285340
X133 2317 2 2312 1 INV1S $T=596440 336120 0 180 $X=595200 $Y=330700
X134 2329 2 2323 1 INV1S $T=597060 315960 0 180 $X=595820 $Y=310540
X135 2337 2 2319 1 INV1S $T=597680 336120 0 180 $X=596440 $Y=330700
X136 2288 2 2339 1 INV1S $T=598300 336120 0 0 $X=598300 $Y=335740
X137 2330 2 2346 1 INV1S $T=602020 326040 0 180 $X=600780 $Y=320620
X138 2354 2 2160 1 INV1S $T=602640 285720 1 180 $X=601400 $Y=285340
X139 2360 2 2331 1 INV1S $T=603260 326040 1 180 $X=602020 $Y=325660
X140 2315 2 2358 1 INV1S $T=602020 336120 0 0 $X=602020 $Y=335740
X141 2355 2 2370 1 INV1S $T=606980 346200 1 0 $X=606980 $Y=340780
X142 2373 2 2366 1 INV1S $T=609460 346200 0 180 $X=608220 $Y=340780
X143 2362 2 2372 1 INV1S $T=608220 346200 0 0 $X=608220 $Y=345820
X144 2376 2 2379 1 INV1S $T=609460 346200 0 0 $X=609460 $Y=345820
X145 2365 2 2385 1 INV1S $T=613180 356280 0 180 $X=611940 $Y=350860
X146 2390 2 2350 1 INV1S $T=613800 336120 1 180 $X=612560 $Y=335740
X147 2363 2 2392 1 INV1S $T=613180 326040 1 0 $X=613180 $Y=320620
X148 2398 2 2417 1 INV1S $T=620000 356280 1 0 $X=620000 $Y=350860
X149 266 2 2419 1 INV1S $T=621240 356280 1 0 $X=621240 $Y=350860
X150 2419 2 422 1 INV1S $T=623720 356280 0 0 $X=623720 $Y=355900
X151 423 2 417 1 INV1S $T=625580 366360 0 180 $X=624340 $Y=360940
X152 423 2 2404 1 INV1S $T=633020 346200 1 180 $X=631780 $Y=345820
X153 423 2 2473 1 INV1S $T=635500 356280 0 0 $X=635500 $Y=355900
X154 2198 2 2432 1 INV1S $T=637360 275640 0 0 $X=637360 $Y=275260
X155 2454 2 2474 1 INV1S $T=637360 326040 1 0 $X=637360 $Y=320620
X156 440 2 2483 1 INV1S $T=644800 275640 1 0 $X=644800 $Y=270220
X157 388 2 2499 1 INV1S $T=646660 305880 0 0 $X=646660 $Y=305500
X158 2499 2 2467 1 INV1S $T=647900 305880 0 0 $X=647900 $Y=305500
X159 440 2 2489 1 INV1S $T=648520 295800 1 0 $X=648520 $Y=290380
X160 440 2 2495 1 INV1S $T=648520 346200 0 0 $X=648520 $Y=345820
X161 440 2 2511 1 INV1S $T=649760 346200 0 0 $X=649760 $Y=345820
X162 2293 2 2521 1 INV1S $T=652240 346200 0 0 $X=652240 $Y=345820
X163 402 2 2526 1 INV1S $T=655960 346200 0 0 $X=655960 $Y=345820
X164 2526 2 2531 1 INV1S $T=657200 356280 1 0 $X=657200 $Y=350860
X165 2499 2 2530 1 INV1S $T=657820 326040 1 0 $X=657820 $Y=320620
X166 461 2 2542 1 INV1S $T=662160 285720 0 0 $X=662160 $Y=285340
X167 460 2 2544 1 INV1S $T=662780 366360 1 0 $X=662780 $Y=360940
X168 2542 2 2547 1 INV1S $T=663400 285720 0 0 $X=663400 $Y=285340
X169 2544 2 464 1 INV1S $T=664020 366360 1 0 $X=664020 $Y=360940
X170 2548 2 2543 1 INV1S $T=665260 285720 1 0 $X=665260 $Y=280300
X171 2614 2 2603 1 INV1S $T=693160 285720 0 180 $X=691920 $Y=280300
X172 2613 2 2617 1 INV1S $T=693160 295800 0 0 $X=693160 $Y=295420
X173 2605 2 2615 1 INV1S $T=693780 275640 0 0 $X=693780 $Y=275260
X174 493 2 2618 1 INV1S $T=698740 305880 0 180 $X=697500 $Y=300460
X175 2622 2 2633 1 INV1S $T=701220 285720 1 0 $X=701220 $Y=280300
X176 501 2 2642 1 INV1S $T=705560 315960 1 180 $X=704320 $Y=315580
X177 2664 2 2640 1 INV1S $T=709280 285720 1 180 $X=708040 $Y=285340
X178 491 2 2654 1 INV1S $T=709900 275640 1 0 $X=709900 $Y=270220
X179 2670 2 2631 1 INV1S $T=711140 305880 1 0 $X=711140 $Y=300460
X180 2682 2 2691 1 INV1S $T=716720 336120 0 0 $X=716720 $Y=335740
X181 2692 2 2663 1 INV1S $T=720440 356280 1 0 $X=720440 $Y=350860
X182 2661 2 2720 1 INV1S $T=724160 326040 1 0 $X=724160 $Y=320620
X183 521 2 2710 1 INV1S $T=727260 275640 1 0 $X=727260 $Y=270220
X184 2698 2 2727 1 INV1S $T=734700 275640 0 0 $X=734700 $Y=275260
X185 2743 2 2705 1 INV1S $T=737800 326040 0 180 $X=736560 $Y=320620
X186 2743 2 498 1 INV1S $T=737800 326040 1 180 $X=736560 $Y=325660
X187 2744 2 2602 1 INV1S $T=738420 295800 1 180 $X=737180 $Y=295420
X188 2735 2 2744 1 INV1S $T=738420 295800 0 0 $X=738420 $Y=295420
X189 2757 2 2731 1 INV1S $T=741520 305880 0 0 $X=741520 $Y=305500
X190 2744 2 2767 1 INV1S $T=743380 295800 0 0 $X=743380 $Y=295420
X191 2795 2 2761 1 INV1S $T=746480 295800 1 180 $X=745240 $Y=295420
X192 2743 2 2773 1 INV1S $T=745240 326040 1 0 $X=745240 $Y=320620
X193 535 2 2781 1 INV1S $T=747100 356280 1 0 $X=747100 $Y=350860
X194 2781 2 2763 1 INV1S $T=750200 346200 0 0 $X=750200 $Y=345820
X195 2781 2 2800 1 INV1S $T=752060 346200 0 0 $X=752060 $Y=345820
X196 2805 2 2772 1 INV1S $T=753920 305880 0 180 $X=752680 $Y=300460
X197 2838 2 2743 1 INV1S $T=767560 315960 1 180 $X=766320 $Y=315580
X198 2845 2 2820 1 INV1S $T=770660 305880 0 0 $X=770660 $Y=305500
X199 2715 2 2838 1 INV1S $T=775620 326040 0 0 $X=775620 $Y=325660
X200 2878 2 2907 1 INV1S $T=789880 346200 0 0 $X=789880 $Y=345820
X201 2903 2 590 1 INV1S $T=792980 265560 1 0 $X=792980 $Y=260140
X202 2914 2 2864 1 INV1S $T=797320 315960 0 0 $X=797320 $Y=315580
X203 2925 2 2872 1 INV1S $T=801040 326040 0 180 $X=799800 $Y=320620
X204 2928 2 2884 1 INV1S $T=801660 336120 1 0 $X=801660 $Y=330700
X205 2898 2 2948 1 INV1S $T=807240 336120 0 0 $X=807240 $Y=335740
X206 617 2 582 1 INV1S $T=812200 366360 0 180 $X=810960 $Y=360940
X207 2963 2 626 1 INV1S $T=819020 265560 0 180 $X=817780 $Y=260140
X208 2960 2 2981 1 INV1S $T=823980 346200 1 0 $X=823980 $Y=340780
X209 2989 2 645 1 INV1S $T=827080 265560 0 180 $X=825840 $Y=260140
X210 2999 2 3001 1 INV1S $T=832660 346200 1 0 $X=832660 $Y=340780
X211 3003 2 3031 1 INV1S $T=851880 346200 1 0 $X=851880 $Y=340780
X212 3060 2 2957 1 INV1S $T=864280 265560 1 180 $X=863040 $Y=265180
X213 3073 2 2993 1 INV1S $T=868620 336120 0 180 $X=867380 $Y=330700
X214 3077 2 3063 1 INV1S $T=870480 336120 0 180 $X=869240 $Y=330700
X215 3073 2 3085 1 INV1S $T=871100 336120 1 0 $X=871100 $Y=330700
X216 3081 2 3072 1 INV1S $T=874820 326040 1 180 $X=873580 $Y=325660
X217 3073 2 3090 1 INV1S $T=878540 315960 1 0 $X=878540 $Y=310540
X218 3082 2 3060 1 INV1S $T=879160 265560 0 0 $X=879160 $Y=265180
X219 3060 2 728 1 INV1S $T=881020 265560 0 0 $X=881020 $Y=265180
X220 3135 2 3119 1 INV1S $T=896520 326040 1 180 $X=895280 $Y=325660
X221 739 2 3136 1 INV1S $T=897760 265560 0 180 $X=896520 $Y=260140
X222 3119 2 3073 1 INV1S $T=896520 326040 0 0 $X=896520 $Y=325660
X223 3073 2 3129 1 INV1S $T=897140 315960 1 0 $X=897140 $Y=310540
X224 741 2 3143 1 INV1S $T=900860 265560 0 180 $X=899620 $Y=260140
X225 3135 2 3125 1 INV1S $T=900240 336120 1 0 $X=900240 $Y=330700
X226 738 2 3135 1 INV1S $T=901480 346200 1 180 $X=900240 $Y=345820
X227 2736 2 3160 1 INV1S $T=907060 275640 0 0 $X=907060 $Y=275260
X228 3160 2 3158 1 INV1S $T=908300 295800 0 180 $X=907060 $Y=290380
X229 3160 2 3180 1 INV1S $T=912020 305880 1 0 $X=912020 $Y=300460
X230 3160 2 752 1 INV1S $T=912640 275640 0 0 $X=912640 $Y=275260
X231 3100 2 3195 1 INV1S $T=921940 346200 0 0 $X=921940 $Y=345820
X232 3125 2 3206 1 INV1S $T=924420 326040 0 0 $X=924420 $Y=325660
X233 3206 2 3197 1 INV1S $T=930000 315960 1 0 $X=930000 $Y=310540
X234 3206 2 3221 1 INV1S $T=930000 315960 0 0 $X=930000 $Y=315580
X235 759 2 3251 1 INV1S $T=944260 356280 0 0 $X=944260 $Y=355900
X236 3251 2 3234 1 INV1S $T=946120 346200 0 0 $X=946120 $Y=345820
X237 3251 2 795 1 INV1S $T=946740 356280 1 0 $X=946740 $Y=350860
X238 819 2 3236 1 INV1S $T=956040 305880 1 180 $X=954800 $Y=305500
X239 819 2 3277 1 INV1S $T=965340 326040 1 0 $X=965340 $Y=320620
X240 786 2 3317 1 INV1S $T=970920 366360 1 0 $X=970920 $Y=360940
X241 3317 2 3286 1 INV1S $T=971540 356280 0 0 $X=971540 $Y=355900
X242 3266 2 3322 1 INV1S $T=975260 285720 1 0 $X=975260 $Y=280300
X243 3277 2 851 1 INV1S $T=975880 346200 0 0 $X=975880 $Y=345820
X244 3235 2 3346 1 INV1S $T=980840 285720 1 0 $X=980840 $Y=280300
X245 3255 2 3351 1 INV1S $T=982080 275640 0 0 $X=982080 $Y=275260
X246 774 2 3366 1 INV1S $T=990140 275640 0 0 $X=990140 $Y=275260
X247 3229 2 892 1 INV1S $T=1000680 275640 1 0 $X=1000680 $Y=270220
X248 803 2 893 1 INV1S $T=1002540 265560 0 180 $X=1001300 $Y=260140
X249 3411 2 3389 1 INV1S $T=1001920 275640 1 0 $X=1001920 $Y=270220
X250 3359 2 877 1 INV1S $T=1003780 285720 0 180 $X=1002540 $Y=280300
X251 851 2 3432 1 INV1S $T=1006260 346200 1 0 $X=1006260 $Y=340780
X252 3350 2 3436 1 INV1S $T=1011840 285720 1 0 $X=1011840 $Y=280300
X253 3189 2 3438 1 INV1S $T=1013080 295800 1 180 $X=1011840 $Y=295420
X254 3227 2 3439 1 INV1S $T=1013700 305880 1 180 $X=1012460 $Y=305500
X255 3409 2 3448 1 INV1S $T=1014320 285720 0 180 $X=1013080 $Y=280300
X256 3420 2 3430 1 INV1S $T=1014940 295800 0 0 $X=1014940 $Y=295420
X257 3264 2 3458 1 INV1S $T=1014940 305880 0 0 $X=1014940 $Y=305500
X258 3281 2 3456 1 INV1S $T=1023620 305880 0 180 $X=1022380 $Y=300460
X259 3482 2 3410 1 INV1S $T=1026100 305880 0 180 $X=1024860 $Y=300460
X260 819 2 3486 1 INV1S $T=1026100 305880 1 0 $X=1026100 $Y=300460
X261 903 2 3504 1 INV1S $T=1031060 356280 1 0 $X=1031060 $Y=350860
X262 3504 2 3510 1 INV1S $T=1032300 356280 1 0 $X=1032300 $Y=350860
X263 939 2 3518 1 INV1S $T=1034780 265560 0 0 $X=1034780 $Y=265180
X264 3504 2 951 1 INV1S $T=1037260 356280 1 0 $X=1037260 $Y=350860
X265 3485 2 3535 1 INV1S $T=1043460 336120 0 0 $X=1043460 $Y=335740
X266 3526 2 3528 1 INV1S $T=1049040 265560 0 0 $X=1049040 $Y=265180
X267 3567 2 3573 1 INV1S $T=1057100 315960 1 0 $X=1057100 $Y=310540
X268 993 2 972 1 INV1S $T=1058960 265560 1 180 $X=1057720 $Y=265180
X269 3535 2 3551 1 INV1S $T=1057720 336120 1 0 $X=1057720 $Y=330700
X270 3535 2 3554 1 INV1S $T=1057720 346200 1 0 $X=1057720 $Y=340780
X271 3560 2 3571 1 INV1S $T=1060200 326040 1 0 $X=1060200 $Y=320620
X272 3592 2 3577 1 INV1S $T=1063300 326040 1 0 $X=1063300 $Y=320620
X273 3602 2 3589 1 INV1S $T=1067020 326040 1 180 $X=1065780 $Y=325660
X274 3568 2 3595 1 INV1S $T=1067020 326040 0 0 $X=1067020 $Y=325660
X275 3530 2 3637 1 INV1S $T=1067640 295800 0 0 $X=1067640 $Y=295420
X276 3616 2 3634 1 INV1S $T=1073840 305880 1 0 $X=1073840 $Y=300460
X277 3622 2 3635 1 INV1S $T=1073840 326040 1 0 $X=1073840 $Y=320620
X278 3630 2 3638 1 INV1S $T=1074460 285720 1 0 $X=1074460 $Y=280300
X279 3639 2 3624 1 INV1S $T=1076940 295800 0 180 $X=1075700 $Y=290380
X280 1008 2 1009 1 INV1S $T=1077560 265560 1 0 $X=1077560 $Y=260140
X281 3650 2 3619 1 INV1S $T=1078800 305880 0 180 $X=1077560 $Y=300460
X282 1013 2 3661 1 INV1S $T=1079420 366360 1 0 $X=1079420 $Y=360940
X283 3663 2 3632 1 INV1S $T=1081280 285720 1 180 $X=1080040 $Y=285340
X284 3598 2 3681 1 INV1S $T=1084380 305880 0 0 $X=1084380 $Y=305500
X285 3666 2 3678 1 INV1S $T=1084380 326040 1 0 $X=1084380 $Y=320620
X286 3667 2 3690 1 INV1S $T=1088100 326040 0 0 $X=1088100 $Y=325660
X287 3691 2 3707 1 INV1S $T=1091820 275640 1 0 $X=1091820 $Y=270220
X288 3714 2 3689 1 INV1S $T=1097400 275640 1 180 $X=1096160 $Y=275260
X289 3637 2 3692 1 INV1S $T=1097400 295800 0 0 $X=1097400 $Y=295420
X290 3723 2 3724 1 INV1S $T=1098640 275640 1 0 $X=1098640 $Y=270220
X291 3637 2 3715 1 INV1S $T=1099880 295800 0 0 $X=1099880 $Y=295420
X292 3730 2 1024 1 INV1S $T=1101740 265560 0 180 $X=1100500 $Y=260140
X293 3730 2 3649 1 INV1S $T=1101740 265560 1 180 $X=1100500 $Y=265180
X294 3732 2 3730 1 INV1S $T=1103600 295800 0 180 $X=1102360 $Y=290380
X295 3749 2 3746 1 INV1S $T=1106080 295800 0 0 $X=1106080 $Y=295420
X296 3756 2 3750 1 INV1S $T=1108560 315960 1 0 $X=1108560 $Y=310540
X297 3748 2 3762 1 INV1S $T=1109180 326040 1 0 $X=1109180 $Y=320620
X298 3720 2 3765 1 INV1S $T=1109800 326040 0 0 $X=1109800 $Y=325660
X299 3753 2 3774 1 INV1S $T=1110420 315960 1 0 $X=1110420 $Y=310540
X300 3761 2 3732 1 INV1S $T=1115380 295800 1 0 $X=1115380 $Y=290380
X301 3739 2 3798 1 INV1S $T=1118480 265560 1 0 $X=1118480 $Y=260140
X302 3779 2 3787 1 INV1S $T=1125300 295800 1 180 $X=1124060 $Y=295420
X303 3802 2 3747 1 INV1S $T=1127780 315960 1 0 $X=1127780 $Y=310540
X304 1055 2 1056 1 INV1S $T=1128400 295800 0 0 $X=1128400 $Y=295420
X305 1055 2 3803 1 INV1S $T=1128400 336120 1 0 $X=1128400 $Y=330700
X306 5 1 2 10 BUF1S $T=220720 285720 1 0 $X=220720 $Y=280300
X307 4 1 2 11 BUF1S $T=220720 305880 1 0 $X=220720 $Y=300460
X308 1109 1 2 1111 BUF1S $T=229400 326040 0 0 $X=229400 $Y=325660
X309 17 1 2 18 BUF1S $T=236220 295800 1 180 $X=233740 $Y=295420
X310 1116 1 2 27 BUF1S $T=235600 265560 0 0 $X=235600 $Y=265180
X311 1094 1 2 1129 BUF1S $T=236220 285720 0 0 $X=236220 $Y=285340
X312 1116 1 2 1132 BUF1S $T=236840 275640 0 0 $X=236840 $Y=275260
X313 25 1 2 1134 BUF1S $T=237460 315960 1 0 $X=237460 $Y=310540
X314 20 1 2 1146 BUF1S $T=240560 346200 0 0 $X=240560 $Y=345820
X315 7 1 2 1149 BUF1S $T=241800 356280 1 0 $X=241800 $Y=350860
X316 31 1 2 1159 BUF1S $T=244280 336120 1 0 $X=244280 $Y=330700
X317 1159 1 2 1154 BUF1S $T=248000 285720 0 180 $X=245520 $Y=280300
X318 39 1 2 36 BUF1S $T=245520 356280 1 0 $X=245520 $Y=350860
X319 1139 1 2 1171 BUF1S $T=247380 315960 0 0 $X=247380 $Y=315580
X320 19 1 2 1173 BUF1S $T=247380 346200 0 0 $X=247380 $Y=345820
X321 1111 1 2 1172 BUF1S $T=249240 326040 1 0 $X=249240 $Y=320620
X322 45 1 2 42 BUF1S $T=249240 356280 1 0 $X=249240 $Y=350860
X323 50 1 2 41 BUF1S $T=254200 346200 1 180 $X=251720 $Y=345820
X324 54 1 2 38 BUF1S $T=258540 356280 0 180 $X=256060 $Y=350860
X325 1129 1 2 1196 BUF1S $T=259780 305880 1 0 $X=259780 $Y=300460
X326 1145 1 2 1217 BUF1S $T=263500 295800 0 0 $X=263500 $Y=295420
X327 1145 1 2 1222 BUF1S $T=265360 315960 1 0 $X=265360 $Y=310540
X328 1216 1 2 1211 BUF1S $T=275900 295800 0 0 $X=275900 $Y=295420
X329 79 1 2 1316 BUF1S $T=305040 326040 0 180 $X=302560 $Y=320620
X330 1316 1 2 95 BUF1S $T=304420 265560 0 0 $X=304420 $Y=265180
X331 100 1 2 1435 BUF1S $T=327360 336120 0 0 $X=327360 $Y=335740
X332 1091 1 2 105 BUF1S $T=333560 305880 1 0 $X=333560 $Y=300460
X333 1435 1 2 108 BUF1S $T=339140 275640 0 0 $X=339140 $Y=275260
X334 103 1 2 1494 BUF1S $T=343480 315960 0 0 $X=343480 $Y=315580
X335 1457 1 2 130 BUF1S $T=347820 275640 0 0 $X=347820 $Y=275260
X336 99 1 2 1515 BUF1S $T=349060 315960 1 0 $X=349060 $Y=310540
X337 1494 1 2 117 BUF1S $T=354020 285720 1 0 $X=354020 $Y=280300
X338 1515 1 2 141 BUF1S $T=358980 265560 0 0 $X=358980 $Y=265180
X339 1524 1 2 1535 BUF1S $T=363320 305880 1 0 $X=363320 $Y=300460
X340 1607 1 2 154 BUF1S $T=383780 295800 1 0 $X=383780 $Y=290380
X341 162 1 2 1653 BUF1S $T=391220 336120 0 0 $X=391220 $Y=335740
X342 160 1 2 1643 BUF1S $T=395560 366360 0 180 $X=393080 $Y=360940
X343 169 1 2 1650 BUF1S $T=394940 346200 0 0 $X=394940 $Y=345820
X344 1655 1 2 1657 BUF1S $T=399280 285720 1 180 $X=396800 $Y=285340
X345 1637 1 2 1632 BUF1S $T=399900 285720 0 0 $X=399900 $Y=285340
X346 180 1 2 1649 BUF1S $T=402380 305880 1 180 $X=399900 $Y=305500
X347 1652 1 2 1624 BUF1S $T=404240 295800 0 180 $X=401760 $Y=290380
X348 179 1 2 1626 BUF1S $T=411680 295800 0 180 $X=409200 $Y=290380
X349 140 1 2 191 BUF1S $T=414160 356280 1 0 $X=414160 $Y=350860
X350 198 1 2 1734 BUF1S $T=422840 356280 1 0 $X=422840 $Y=350860
X351 144 1 2 204 BUF1S $T=426560 315960 1 0 $X=426560 $Y=310540
X352 211 1 2 212 BUF1S $T=428420 326040 0 0 $X=428420 $Y=325660
X353 194 1 2 215 BUF1S $T=430900 295800 0 0 $X=430900 $Y=295420
X354 227 1 2 224 BUF1S $T=447020 265560 0 180 $X=444540 $Y=260140
X355 199 1 2 1796 BUF1S $T=446400 326040 0 0 $X=446400 $Y=325660
X356 208 1 2 1806 BUF1S $T=447020 265560 1 0 $X=447020 $Y=260140
X357 234 1 2 1808 BUF1S $T=447640 356280 0 0 $X=447640 $Y=355900
X358 223 1 2 1864 BUF1S $T=453220 305880 1 0 $X=453220 $Y=300460
X359 230 1 2 1835 BUF1S $T=455080 346200 0 0 $X=455080 $Y=345820
X360 195 1 2 241 BUF1S $T=456940 295800 1 0 $X=456940 $Y=290380
X361 1734 1 2 251 BUF1S $T=467480 275640 0 0 $X=467480 $Y=275260
X362 260 1 2 1901 BUF1S $T=477400 346200 1 0 $X=477400 $Y=340780
X363 246 1 2 274 BUF1S $T=492280 295800 1 0 $X=492280 $Y=290380
X364 204 1 2 279 BUF1S $T=495380 315960 0 0 $X=495380 $Y=315580
X365 1868 1 2 285 BUF1S $T=496000 305880 1 0 $X=496000 $Y=300460
X366 1901 1 2 1987 BUF1S $T=506540 305880 1 0 $X=506540 $Y=300460
X367 1779 1 2 2000 BUF1S $T=510260 275640 1 0 $X=510260 $Y=270220
X368 1886 1 2 292 BUF1S $T=511500 295800 1 0 $X=511500 $Y=290380
X369 140 1 2 2040 BUF1S $T=518940 356280 0 0 $X=518940 $Y=355900
X370 2074 1 2 1989 BUF1S $T=530720 336120 0 180 $X=528240 $Y=330700
X371 2089 1 2 2012 BUF1S $T=530720 336120 1 180 $X=528240 $Y=335740
X372 2115 1 2 2025 BUF1S $T=540640 346200 1 180 $X=538160 $Y=345820
X373 2133 1 2 2095 BUF1S $T=544360 356280 0 180 $X=541880 $Y=350860
X374 2162 1 2 2089 BUF1S $T=549320 336120 0 0 $X=549320 $Y=335740
X375 2169 1 2 2074 BUF1S $T=551180 336120 1 0 $X=551180 $Y=330700
X376 2180 1 2 2115 BUF1S $T=555520 346200 0 180 $X=553040 $Y=340780
X377 212 1 2 2185 BUF1S $T=554280 326040 0 0 $X=554280 $Y=325660
X378 1796 1 2 2208 BUF1S $T=556760 326040 0 0 $X=556760 $Y=325660
X379 2133 1 2 2200 BUF1S $T=562340 356280 0 180 $X=559860 $Y=350860
X380 2216 1 2 2162 BUF1S $T=564200 336120 0 180 $X=561720 $Y=330700
X381 356 1 2 2133 BUF1S $T=566060 366360 0 180 $X=563580 $Y=360940
X382 363 1 2 2180 BUF1S $T=571020 346200 1 180 $X=568540 $Y=345820
X383 369 1 2 2216 BUF1S $T=571020 356280 0 0 $X=571020 $Y=355900
X384 367 1 2 2169 BUF1S $T=574120 336120 0 0 $X=574120 $Y=335740
X385 2251 1 2 2257 BUF1S $T=579080 275640 0 0 $X=579080 $Y=275260
X386 388 1 2 2202 BUF1S $T=585280 275640 0 0 $X=585280 $Y=275260
X387 1808 1 2 391 BUF1S $T=587760 275640 0 0 $X=587760 $Y=275260
X388 2270 1 2 396 BUF1S $T=590240 295800 0 0 $X=590240 $Y=295420
X389 2185 1 2 425 BUF1S $T=625580 366360 1 0 $X=625580 $Y=360940
X390 241 1 2 427 BUF1S $T=631160 295800 1 0 $X=631160 $Y=290380
X391 194 1 2 428 BUF1S $T=631160 366360 1 0 $X=631160 $Y=360940
X392 2239 1 2 2445 BUF1S $T=633020 315960 0 0 $X=633020 $Y=315580
X393 1835 1 2 2470 BUF1S $T=635500 285720 0 0 $X=635500 $Y=285340
X394 1864 1 2 436 BUF1S $T=636740 275640 1 0 $X=636740 $Y=270220
X395 2040 1 2 421 BUF1S $T=645420 356280 0 0 $X=645420 $Y=355900
X396 470 1 2 476 BUF1S $T=682620 356280 0 0 $X=682620 $Y=355900
X397 491 1 2 503 BUF1S $T=709900 265560 0 180 $X=707420 $Y=260140
X398 2675 1 2 483 BUF1S $T=711760 275640 1 180 $X=709280 $Y=275260
X399 2683 1 2 2653 BUF1S $T=714240 336120 0 0 $X=714240 $Y=335740
X400 2686 1 2 2677 BUF1S $T=716100 326040 1 0 $X=716100 $Y=320620
X401 513 1 2 509 BUF1S $T=718580 265560 1 0 $X=718580 $Y=260140
X402 2702 1 2 2684 BUF1S $T=719820 265560 0 0 $X=719820 $Y=265180
X403 2678 1 2 2675 BUF1S $T=722300 326040 0 180 $X=719820 $Y=320620
X404 2704 1 2 2701 BUF1S $T=722920 275640 1 0 $X=722920 $Y=270220
X405 520 1 2 2678 BUF1S $T=725400 356280 0 180 $X=722920 $Y=350860
X406 2678 1 2 522 BUF1S $T=725400 356280 1 0 $X=725400 $Y=350860
X407 522 1 2 2735 BUF1S $T=734080 346200 0 0 $X=734080 $Y=345820
X408 2602 1 2 526 BUF1S $T=738420 275640 0 180 $X=735940 $Y=270220
X409 2746 1 2 2738 BUF1S $T=738420 305880 1 0 $X=738420 $Y=300460
X410 2751 1 2 2698 BUF1S $T=739660 285720 1 0 $X=739660 $Y=280300
X411 518 1 2 2765 BUF1S $T=740900 326040 1 0 $X=740900 $Y=320620
X412 539 1 2 2780 BUF1S $T=746480 346200 0 0 $X=746480 $Y=345820
X413 558 1 2 559 BUF1S $T=759500 366360 1 0 $X=759500 $Y=360940
X414 2821 1 2 2818 BUF1S $T=761360 356280 1 0 $X=761360 $Y=350860
X415 2793 1 2 2810 BUF1S $T=765080 356280 1 180 $X=762600 $Y=355900
X416 2767 1 2 2833 BUF1S $T=769420 295800 1 0 $X=769420 $Y=290380
X417 582 1 2 2793 BUF1S $T=786160 346200 1 180 $X=783680 $Y=345820
X418 2762 1 2 2882 BUF1S $T=789880 305880 0 0 $X=789880 $Y=305500
X419 2942 1 2 2623 BUF1S $T=817160 315960 1 180 $X=814680 $Y=315580
X420 2882 1 2 2971 BUF1S $T=819640 315960 1 0 $X=819640 $Y=310540
X421 2993 1 2 2909 BUF1S $T=837000 326040 0 180 $X=834520 $Y=320620
X422 2971 1 2 3014 BUF1S $T=837000 315960 1 0 $X=837000 $Y=310540
X423 2942 1 2 3004 BUF1S $T=837000 326040 1 0 $X=837000 $Y=320620
X424 2993 1 2 2915 BUF1S $T=840720 326040 1 0 $X=840720 $Y=320620
X425 3045 1 2 3030 BUF1S $T=856220 326040 1 0 $X=856220 $Y=320620
X426 717 1 2 2911 BUF1S $T=876680 265560 1 180 $X=874200 $Y=265180
X427 3090 1 2 3024 BUF1S $T=876680 305880 1 180 $X=874200 $Y=305500
X428 3014 1 2 3099 BUF1S $T=877920 295800 0 0 $X=877920 $Y=295420
X429 723 1 2 3041 BUF1S $T=880400 356280 0 180 $X=877920 $Y=350860
X430 726 1 2 3044 BUF1S $T=890940 346200 0 0 $X=890940 $Y=345820
X431 3137 1 2 3061 BUF1S $T=899000 285720 0 180 $X=896520 $Y=280300
X432 740 1 2 738 BUF1S $T=899620 356280 1 180 $X=897140 $Y=355900
X433 710 1 2 3145 BUF1S $T=897760 346200 0 0 $X=897760 $Y=345820
X434 3138 1 2 3151 BUF1S $T=901480 315960 0 0 $X=901480 $Y=315580
X435 3137 1 2 744 BUF1S $T=908300 275640 1 0 $X=908300 $Y=270220
X436 3173 1 2 3164 BUF1S $T=910780 305880 0 0 $X=910780 $Y=305500
X437 3178 1 2 3126 BUF1S $T=911400 315960 0 0 $X=911400 $Y=315580
X438 3180 1 2 3174 BUF1S $T=915120 326040 0 0 $X=915120 $Y=325660
X439 3176 1 2 3171 BUF1S $T=915740 315960 1 0 $X=915740 $Y=310540
X440 724 1 2 3203 BUF1S $T=921940 356280 0 0 $X=921940 $Y=355900
X441 3209 1 2 3137 BUF1S $T=926280 285720 0 180 $X=923800 $Y=280300
X442 3227 1 2 3215 BUF1S $T=932480 315960 1 0 $X=932480 $Y=310540
X443 3209 1 2 766 BUF1S $T=933100 265560 0 0 $X=933100 $Y=265180
X444 3189 1 2 3242 BUF1S $T=934960 305880 0 0 $X=934960 $Y=305500
X445 2747 1 2 791 BUF1S $T=936200 275640 0 0 $X=936200 $Y=275260
X446 792 1 2 3237 BUF1S $T=940540 285720 1 180 $X=938060 $Y=285340
X447 3236 1 2 3209 BUF1S $T=941160 295800 1 180 $X=938680 $Y=295420
X448 726 1 2 806 BUF1S $T=947980 346200 0 0 $X=947980 $Y=345820
X449 3254 1 2 3218 BUF1S $T=951080 305880 1 180 $X=948600 $Y=305500
X450 791 1 2 3253 BUF1S $T=949220 275640 0 0 $X=949220 $Y=275260
X451 3253 1 2 3254 BUF1S $T=953560 305880 1 180 $X=951080 $Y=305500
X452 3145 1 2 3291 BUF1S $T=966580 346200 0 0 $X=966580 $Y=345820
X453 3409 1 2 846 BUF1S $T=1001300 275640 1 180 $X=998820 $Y=275260
X454 877 1 2 3396 BUF1S $T=1001920 285720 0 0 $X=1001920 $Y=285340
X455 3420 1 2 840 BUF1S $T=1005020 265560 1 180 $X=1002540 $Y=265180
X456 3389 1 2 3368 BUF1S $T=1002540 275640 0 0 $X=1002540 $Y=275260
X457 3410 1 2 882 BUF1S $T=1006260 285720 0 180 $X=1003780 $Y=280300
X458 3436 1 2 3354 BUF1S $T=1008740 285720 0 180 $X=1006260 $Y=280300
X459 910 1 2 3350 BUF1S $T=1013700 265560 0 180 $X=1011220 $Y=260140
X460 913 1 2 3369 BUF1S $T=1016180 356280 0 0 $X=1016180 $Y=355900
X461 925 1 2 902 BUF1S $T=1026100 366360 0 180 $X=1023620 $Y=360940
X462 3432 1 2 3485 BUF1S $T=1025480 346200 1 0 $X=1025480 $Y=340780
X463 3486 1 2 915 BUF1S $T=1027340 285720 1 0 $X=1027340 $Y=280300
X464 939 1 2 934 BUF1S $T=1031680 265560 1 180 $X=1029200 $Y=265180
X465 944 1 2 3506 BUF1S $T=1034780 265560 1 180 $X=1032300 $Y=265180
X466 945 1 2 881 BUF1S $T=1034780 366360 0 180 $X=1032300 $Y=360940
X467 3518 1 2 958 BUF1S $T=1039740 265560 1 0 $X=1039740 $Y=260140
X468 3485 1 2 943 BUF1S $T=1042220 356280 0 0 $X=1042220 $Y=355900
X469 3537 1 2 964 BUF1S $T=1045940 275640 1 180 $X=1043460 $Y=275260
X470 3486 1 2 3530 BUF1S $T=1043460 295800 0 0 $X=1043460 $Y=295420
X471 3526 1 2 970 BUF1S $T=1048420 275640 0 180 $X=1045940 $Y=270220
X472 3530 1 2 3529 BUF1S $T=1046560 295800 0 0 $X=1046560 $Y=295420
X473 3548 1 2 3526 BUF1S $T=1052760 275640 1 180 $X=1050280 $Y=275260
X474 3531 1 2 975 BUF1S $T=1050280 285720 0 0 $X=1050280 $Y=285340
X475 3581 1 2 3521 BUF1S $T=1060820 275640 1 0 $X=1060820 $Y=270220
X476 3581 1 2 993 BUF1S $T=1066400 275640 0 180 $X=1063920 $Y=270220
X477 3611 1 2 983 BUF1S $T=1068880 265560 1 180 $X=1066400 $Y=265180
X478 3612 1 2 3584 BUF1S $T=1069500 336120 0 0 $X=1069500 $Y=335740
X479 3484 1 2 3636 BUF1S $T=1072600 315960 1 0 $X=1072600 $Y=310540
X480 3484 1 2 3596 BUF1S $T=1073220 315960 0 0 $X=1073220 $Y=315580
X481 1007 1 2 932 BUF1S $T=1077560 265560 0 180 $X=1075080 $Y=260140
X482 1011 1 2 3549 BUF1S $T=1079420 366360 0 180 $X=1076940 $Y=360940
X483 3649 1 2 3547 BUF1S $T=1084380 275640 1 180 $X=1081900 $Y=275260
X484 3607 1 2 3655 BUF1S $T=1086240 295800 0 180 $X=1083760 $Y=290380
X485 3529 1 2 1019 BUF1S $T=1088100 265560 0 180 $X=1085620 $Y=260140
X486 3551 1 2 3721 BUF1S $T=1098020 336120 0 0 $X=1098020 $Y=335740
X487 3725 1 2 3726 BUF1S $T=1098640 285720 0 0 $X=1098640 $Y=285340
X488 3716 1 2 3722 BUF1S $T=1099880 295800 1 0 $X=1099880 $Y=290380
X489 3732 1 2 3627 BUF1S $T=1107320 326040 0 0 $X=1107320 $Y=325660
X490 3636 1 2 3761 BUF1S $T=1107940 295800 1 0 $X=1107940 $Y=290380
X491 3721 1 2 3737 BUF1S $T=1114140 346200 0 0 $X=1114140 $Y=345820
X492 3761 1 2 1040 BUF1S $T=1118480 265560 1 180 $X=1116000 $Y=265180
X493 3783 1 2 3791 BUF1S $T=1119100 326040 0 0 $X=1119100 $Y=325660
X494 3715 1 2 1038 BUF1S $T=1126540 285720 1 0 $X=1126540 $Y=280300
X495 3801 1 2 3797 BUF1S $T=1127160 265560 0 0 $X=1127160 $Y=265180
X496 1082 1 2 1085 DELB $T=223820 346200 1 0 $X=223820 $Y=340780
X497 1087 1 2 1077 DELB $T=224440 275640 0 0 $X=224440 $Y=275260
X498 1108 1 2 1096 DELB $T=231260 305880 1 0 $X=231260 $Y=300460
X499 1487 1 2 1492 DELB $T=344720 295800 1 0 $X=344720 $Y=290380
X500 2572 1 2 2580 DELB $T=675800 275640 1 0 $X=675800 $Y=270220
X501 479 1 2 481 DELB $T=680140 265560 1 0 $X=680140 $Y=260140
X502 2604 1 2 2587 DELB $T=688200 265560 1 0 $X=688200 $Y=260140
X503 2616 1 2 2619 DELB $T=694400 295800 1 0 $X=694400 $Y=290380
X504 2621 1 2 2637 DELB $T=698740 265560 1 0 $X=698740 $Y=260140
X505 2672 1 2 2682 DELB $T=709280 336120 0 0 $X=709280 $Y=335740
X506 2679 1 2 2693 DELB $T=713000 305880 0 0 $X=713000 $Y=305500
X507 504 1 2 517 DELB $T=717340 356280 0 0 $X=717340 $Y=355900
X508 530 1 2 536 DELB $T=737180 356280 1 0 $X=737180 $Y=350860
X509 2755 1 2 2749 DELB $T=742760 326040 0 0 $X=742760 $Y=325660
X510 543 1 2 545 DELB $T=747720 336120 0 0 $X=747720 $Y=335740
X511 552 1 2 562 DELB $T=757640 336120 0 0 $X=757640 $Y=335740
X512 546 1 2 568 DELB $T=765700 336120 0 0 $X=765700 $Y=335740
X513 2854 1 2 2853 DELB $T=774380 305880 0 0 $X=774380 $Y=305500
X514 575 1 2 2868 DELB $T=777480 336120 0 0 $X=777480 $Y=335740
X515 2860 1 2 2840 DELB $T=778100 315960 1 0 $X=778100 $Y=310540
X516 578 1 2 2887 DELB $T=779960 356280 0 0 $X=779960 $Y=355900
X517 2886 1 2 2898 DELB $T=784300 336120 1 0 $X=784300 $Y=330700
X518 2888 1 2 2892 DELB $T=786160 295800 0 0 $X=786160 $Y=295420
X519 588 1 2 594 DELB $T=791120 326040 0 0 $X=791120 $Y=325660
X520 2919 1 2 2936 DELB $T=798560 315960 1 0 $X=798560 $Y=310540
X521 2910 1 2 2933 DELB $T=801040 326040 0 0 $X=801040 $Y=325660
X522 2940 1 2 2941 DELB $T=804140 305880 0 0 $X=804140 $Y=305500
X523 2951 1 2 2956 DELB $T=810960 305880 0 0 $X=810960 $Y=305500
X524 2961 1 2 2960 DELB $T=817780 356280 0 0 $X=817780 $Y=355900
X525 2977 1 2 2978 DELB $T=823360 295800 0 0 $X=823360 $Y=295420
X526 639 1 2 647 DELB $T=823360 336120 1 0 $X=823360 $Y=330700
X527 644 1 2 655 DELB $T=828320 356280 0 0 $X=828320 $Y=355900
X528 2997 1 2 3010 DELB $T=832040 315960 1 0 $X=832040 $Y=310540
X529 2996 1 2 3009 DELB $T=832660 295800 0 0 $X=832660 $Y=295420
X530 3005 1 2 2999 DELB $T=834520 356280 1 0 $X=834520 $Y=350860
X531 670 1 2 676 DELB $T=840100 326040 0 0 $X=840100 $Y=325660
X532 677 1 2 684 DELB $T=845680 326040 0 0 $X=845680 $Y=325660
X533 681 1 2 692 DELB $T=849400 336120 1 0 $X=849400 $Y=330700
X534 3025 1 2 3036 DELB $T=850020 295800 0 0 $X=850020 $Y=295420
X535 3092 1 2 3094 DELB $T=876060 336120 1 0 $X=876060 $Y=330700
X536 3107 1 2 3106 DELB $T=881020 285720 0 0 $X=881020 $Y=285340
X537 3102 1 2 3111 DELB $T=885360 295800 0 0 $X=885360 $Y=295420
X538 3110 1 2 3131 DELB $T=890940 285720 0 0 $X=890940 $Y=285340
X539 3120 1 2 3130 DELB $T=892180 315960 1 0 $X=892180 $Y=310540
X540 3133 1 2 3132 DELB $T=895280 336120 1 0 $X=895280 $Y=330700
X541 3128 1 2 3148 DELB $T=900240 295800 1 0 $X=900240 $Y=290380
X542 747 1 2 749 DELB $T=905820 295800 0 0 $X=905820 $Y=295420
X543 746 1 2 3150 DELB $T=906440 336120 1 0 $X=906440 $Y=330700
X544 3140 1 2 3156 DELB $T=909540 336120 0 0 $X=909540 $Y=335740
X545 3172 1 2 755 DELB $T=910160 265560 0 0 $X=910160 $Y=265180
X546 756 1 2 763 DELB $T=915740 295800 0 0 $X=915740 $Y=295420
X547 3184 1 2 3185 DELB $T=916980 336120 0 0 $X=916980 $Y=335740
X548 767 1 2 775 DELB $T=923800 366360 1 0 $X=923800 $Y=360940
X549 753 1 2 3187 DELB $T=926280 305880 0 0 $X=926280 $Y=305500
X550 776 1 2 784 DELB $T=930000 366360 1 0 $X=930000 $Y=360940
X551 3233 1 2 3194 DELB $T=934960 295800 1 0 $X=934960 $Y=290380
X552 3240 1 2 3222 DELB $T=937440 326040 0 0 $X=937440 $Y=325660
X553 798 1 2 805 DELB $T=945500 326040 1 0 $X=945500 $Y=320620
X554 799 1 2 813 DELB $T=947360 356280 0 0 $X=947360 $Y=355900
X555 3259 1 2 3271 DELB $T=949840 356280 1 0 $X=949840 $Y=350860
X556 810 1 2 820 DELB $T=951700 315960 1 0 $X=951700 $Y=310540
X557 827 1 2 831 DELB $T=961000 336120 1 0 $X=961000 $Y=330700
X558 3273 1 2 3298 DELB $T=965340 346200 1 0 $X=965340 $Y=340780
X559 832 1 2 841 DELB $T=965340 366360 1 0 $X=965340 $Y=360940
X560 3269 1 2 3315 DELB $T=970920 346200 1 0 $X=970920 $Y=340780
X561 847 1 2 3319 DELB $T=974020 356280 0 0 $X=974020 $Y=355900
X562 814 1 2 3313 DELB $T=977120 346200 0 0 $X=977120 $Y=345820
X563 856 1 2 861 DELB $T=980220 336120 0 0 $X=980220 $Y=335740
X564 860 1 2 867 DELB $T=981460 326040 1 0 $X=981460 $Y=320620
X565 872 1 2 880 DELB $T=987660 346200 0 0 $X=987660 $Y=345820
X566 3362 1 2 3384 DELB $T=989520 356280 0 0 $X=989520 $Y=355900
X567 895 1 2 3424 DELB $T=1002540 356280 1 0 $X=1002540 $Y=350860
X568 3383 1 2 3413 DELB $T=1006880 346200 0 0 $X=1006880 $Y=345820
X569 3475 1 2 3476 DELB $T=1021760 356280 1 0 $X=1021760 $Y=350860
X570 937 1 2 955 DELB $T=1036020 366360 1 0 $X=1036020 $Y=360940
X571 948 1 2 966 DELB $T=1039740 346200 0 0 $X=1039740 $Y=345820
X572 960 1 2 973 DELB $T=1042220 315960 0 0 $X=1042220 $Y=315580
X573 3531 1 2 3543 DELB $T=1043460 285720 0 0 $X=1043460 $Y=285340
X574 971 1 2 981 DELB $T=1047800 366360 1 0 $X=1047800 $Y=360940
X575 3545 1 2 3544 DELB $T=1048420 315960 1 0 $X=1048420 $Y=310540
X576 3550 1 2 3558 DELB $T=1050900 315960 0 0 $X=1050900 $Y=315580
X577 979 1 2 3562 DELB $T=1050900 326040 0 0 $X=1050900 $Y=325660
X578 3561 1 2 3575 DELB $T=1058960 366360 1 0 $X=1058960 $Y=360940
X579 994 1 2 998 DELB $T=1062680 346200 1 0 $X=1062680 $Y=340780
X580 3557 1 2 3574 DELB $T=1063300 356280 0 0 $X=1063300 $Y=355900
X581 997 1 2 1001 DELB $T=1066400 346200 0 0 $X=1066400 $Y=345820
X582 996 1 2 1006 DELB $T=1070120 356280 0 0 $X=1070120 $Y=355900
X583 3606 1 2 3640 DELB $T=1075080 346200 0 0 $X=1075080 $Y=345820
X584 3658 1 2 3675 DELB $T=1079420 326040 1 0 $X=1079420 $Y=320620
X585 3683 1 2 3691 DELB $T=1086860 285720 1 0 $X=1086860 $Y=280300
X586 3693 1 2 3709 DELB $T=1089960 356280 0 0 $X=1089960 $Y=355900
X587 3711 1 2 3713 DELB $T=1094920 326040 1 0 $X=1094920 $Y=320620
X588 3660 1 2 3704 DELB $T=1094920 346200 1 0 $X=1094920 $Y=340780
X589 1033 1 2 1039 DELB $T=1107940 346200 0 0 $X=1107940 $Y=345820
X590 3771 1 2 1034 DELB $T=1111660 275640 1 0 $X=1111660 $Y=270220
X591 3768 1 2 3780 DELB $T=1111660 366360 1 0 $X=1111660 $Y=360940
X592 3744 1 2 3698 DELB $T=1116000 336120 1 0 $X=1116000 $Y=330700
X593 3777 1 2 3800 DELB $T=1116620 295800 1 0 $X=1116620 $Y=290380
X594 1045 1 2 1049 DELB $T=1116620 346200 0 0 $X=1116620 $Y=345820
X595 3792 1 2 3790 DELB $T=1117240 285720 1 0 $X=1117240 $Y=280300
X596 1083 1 2 1092 DELA $T=224440 305880 0 0 $X=224440 $Y=305500
X597 1409 1 2 1431 DELA $T=324880 336120 1 0 $X=324880 $Y=330700
X598 1420 1 2 1406 DELA $T=325500 356280 0 0 $X=325500 $Y=355900
X599 1448 1 2 1460 DELA $T=331700 295800 0 0 $X=331700 $Y=295420
X600 1462 1 2 1455 DELA $T=336040 326040 0 0 $X=336040 $Y=325660
X601 1436 1 2 1432 DELA $T=342860 356280 1 0 $X=342860 $Y=350860
X602 125 1 2 1483 DELA $T=356500 275640 1 0 $X=356500 $Y=270220
X603 1529 1 2 1542 DELA $T=357740 295800 0 0 $X=357740 $Y=295420
X604 190 1 2 1697 DELA $T=414780 265560 0 0 $X=414780 $Y=265180
X605 2649 1 2 2674 DELA $T=706180 315960 0 0 $X=706180 $Y=315580
X606 2658 1 2 2624 DELA $T=709280 265560 0 0 $X=709280 $Y=265180
X607 510 1 2 514 DELA $T=714240 346200 0 0 $X=714240 $Y=345820
X608 2688 1 2 2700 DELA $T=716720 315960 0 0 $X=716720 $Y=315580
X609 2697 1 2 2711 DELA $T=718580 305880 0 0 $X=718580 $Y=305500
X610 2704 1 2 2702 DELA $T=721060 295800 1 0 $X=721060 $Y=290380
X611 525 1 2 528 DELA $T=729120 356280 1 0 $X=729120 $Y=350860
X612 2740 1 2 2745 DELA $T=737800 326040 0 0 $X=737800 $Y=325660
X613 538 1 2 541 DELA $T=742140 356280 1 0 $X=742140 $Y=350860
X614 2776 1 2 2791 DELA $T=746480 326040 1 0 $X=746480 $Y=320620
X615 2798 1 2 2786 DELA $T=752680 336120 0 0 $X=752680 $Y=335740
X616 2834 1 2 2841 DELA $T=765700 305880 0 0 $X=765700 $Y=305500
X617 595 1 2 602 DELA $T=796080 326040 0 0 $X=796080 $Y=325660
X618 2973 1 2 2975 DELA $T=826460 315960 1 0 $X=826460 $Y=310540
X619 658 1 2 667 DELA $T=835140 326040 0 0 $X=835140 $Y=325660
X620 664 1 2 673 DELA $T=837620 295800 0 0 $X=837620 $Y=295420
X621 3020 1 2 3027 DELA $T=845680 305880 1 0 $X=845680 $Y=300460
X622 3087 1 2 3097 DELA $T=873580 285720 1 0 $X=873580 $Y=280300
X623 3093 1 2 3101 DELA $T=876060 285720 0 0 $X=876060 $Y=285340
X624 3118 1 2 3123 DELA $T=885980 285720 0 0 $X=885980 $Y=285340
X625 734 1 2 736 DELA $T=892800 305880 0 0 $X=892800 $Y=305500
X626 3134 1 2 3144 DELA $T=895280 295800 1 0 $X=895280 $Y=290380
X627 3139 1 2 3155 DELA $T=901480 336120 1 0 $X=901480 $Y=330700
X628 745 1 2 748 DELA $T=904580 326040 1 0 $X=904580 $Y=320620
X629 3235 1 2 3224 DELA $T=935580 265560 0 0 $X=935580 $Y=265180
X630 789 1 2 794 DELA $T=937440 356280 1 0 $X=937440 $Y=350860
X631 797 1 2 802 DELA $T=944260 265560 0 0 $X=944260 $Y=265180
X632 3255 1 2 3256 DELA $T=947360 275640 1 0 $X=947360 $Y=270220
X633 3266 1 2 3258 DELA $T=951700 275640 0 0 $X=951700 $Y=275260
X634 811 1 2 826 DELA $T=956040 336120 1 0 $X=956040 $Y=330700
X635 3281 1 2 3267 DELA $T=960380 275640 0 0 $X=960380 $Y=275260
X636 3264 1 2 3257 DELA $T=964100 275640 1 0 $X=964100 $Y=270220
X637 3349 1 2 3353 DELA $T=982700 346200 0 0 $X=982700 $Y=345820
X638 864 1 2 874 DELA $T=985180 336120 0 0 $X=985180 $Y=335740
X639 870 1 2 878 DELA $T=987040 326040 1 0 $X=987040 $Y=320620
X640 884 1 2 891 DELA $T=993860 356280 1 0 $X=993860 $Y=350860
X641 886 1 2 894 DELA $T=996340 346200 0 0 $X=996340 $Y=345820
X642 889 1 2 897 DELA $T=996960 295800 0 0 $X=996960 $Y=295420
X643 3421 1 2 3440 DELA $T=1004400 336120 0 0 $X=1004400 $Y=335740
X644 900 1 2 907 DELA $T=1005640 326040 1 0 $X=1005640 $Y=320620
X645 909 1 2 3459 DELA $T=1015560 346200 0 0 $X=1015560 $Y=345820
X646 918 1 2 924 DELA $T=1020520 346200 1 0 $X=1020520 $Y=340780
X647 3491 1 2 3514 DELA $T=1031060 315960 0 0 $X=1031060 $Y=315580
X648 950 1 2 959 DELA $T=1037880 315960 1 0 $X=1037880 $Y=310540
X649 957 1 2 974 DELA $T=1040980 366360 1 0 $X=1040980 $Y=360940
X650 3537 1 2 3541 DELA $T=1045320 285720 1 0 $X=1045320 $Y=280300
X651 3548 1 2 3570 DELA $T=1052760 285720 0 0 $X=1052760 $Y=285340
X652 3580 1 2 3572 DELA $T=1064540 326040 1 0 $X=1064540 $Y=320620
X653 3641 1 2 3654 DELA $T=1078800 295800 0 0 $X=1078800 $Y=295420
X654 3682 1 2 3697 DELA $T=1086860 275640 1 0 $X=1086860 $Y=270220
X655 3674 1 2 3668 DELA $T=1089960 326040 1 0 $X=1089960 $Y=320620
X656 3684 1 2 3688 DELA $T=1090580 315960 1 0 $X=1090580 $Y=310540
X657 1037 1 2 1042 DELA $T=1110420 336120 0 0 $X=1110420 $Y=335740
X658 3767 1 2 3782 DELA $T=1111040 305880 0 0 $X=1111040 $Y=305500
X659 3784 1 2 3785 DELA $T=1120960 336120 1 0 $X=1120960 $Y=330700
X660 1050 1 2 1053 DELA $T=1121580 346200 0 0 $X=1121580 $Y=345820
X661 1076 8 17 2 1 1072 QDFFRBN $T=220720 326040 1 0 $X=220720 $Y=320620
X662 1078 8 18 2 1 21 QDFFRBN $T=221340 265560 1 0 $X=221340 $Y=260140
X663 1079 8 18 2 1 1073 QDFFRBN $T=221340 275640 1 0 $X=221340 $Y=270220
X664 1074 8 18 2 1 1094 QDFFRBN $T=221340 295800 1 0 $X=221340 $Y=290380
X665 1080 8 17 2 1 1107 QDFFRBN $T=221340 315960 1 0 $X=221340 $Y=310540
X666 1081 8 17 2 1 1075 QDFFRBN $T=221340 336120 0 0 $X=221340 $Y=335740
X667 1385 8 103 2 1 1436 QDFFRBN $T=318680 346200 0 0 $X=318680 $Y=345820
X668 1414 8 103 2 1 1420 QDFFRBN $T=324260 366360 1 0 $X=324260 $Y=360940
X669 1438 8 103 2 1 1409 QDFFRBN $T=329220 346200 1 0 $X=329220 $Y=340780
X670 1454 8 103 2 1 1462 QDFFRBN $T=333560 336120 1 0 $X=333560 $Y=330700
X671 1465 8 1494 2 1 1448 QDFFRBN $T=336040 305880 1 0 $X=336040 $Y=300460
X672 1466 8 103 2 1 1484 QDFFRBN $T=336040 326040 1 0 $X=336040 $Y=320620
X673 1468 8 1494 2 1 1464 QDFFRBN $T=337280 305880 0 0 $X=337280 $Y=305500
X674 109 8 117 2 1 121 QDFFRBN $T=339140 265560 1 0 $X=339140 $Y=260140
X675 1493 8 1494 2 1 1487 QDFFRBN $T=354020 295800 1 180 $X=342240 $Y=295420
X676 1495 8 117 2 1 125 QDFFRBN $T=344720 275640 1 0 $X=344720 $Y=270220
X677 1500 8 1494 2 1 1524 QDFFRBN $T=347820 305880 1 0 $X=347820 $Y=300460
X678 1542 8 1494 2 1 1512 QDFFRBN $T=363320 285720 1 180 $X=351540 $Y=285340
X679 1510 8 117 2 1 1504 QDFFRBN $T=368280 275640 1 180 $X=356500 $Y=275260
X680 1955 280 286 2 1 288 QDFFRBN $T=497240 366360 1 0 $X=497240 $Y=360940
X681 297 280 286 2 1 289 QDFFRBN $T=521420 366360 0 180 $X=509640 $Y=360940
X682 2578 480 2602 2 1 2604 QDFFRBN $T=679520 265560 0 0 $X=679520 $Y=265180
X683 2580 480 2602 2 1 2592 QDFFRBN $T=679520 285720 1 0 $X=679520 $Y=280300
X684 2619 480 2602 2 1 2600 QDFFRBN $T=698740 285720 1 180 $X=686960 $Y=285340
X685 2624 480 483 2 1 482 QDFFRBN $T=700600 275640 0 180 $X=688820 $Y=270220
X686 2643 480 2675 2 1 2686 QDFFRBN $T=704320 326040 1 0 $X=704320 $Y=320620
X687 2644 480 2678 2 1 2685 QDFFRBN $T=704320 336120 1 0 $X=704320 $Y=330700
X688 2645 480 2678 2 1 2672 QDFFRBN $T=704320 346200 1 0 $X=704320 $Y=340780
X689 2657 480 2678 2 1 2692 QDFFRBN $T=706180 356280 1 0 $X=706180 $Y=350860
X690 2674 480 2675 2 1 501 QDFFRBN $T=719820 315960 0 180 $X=708040 $Y=310540
X691 515 480 508 2 1 504 QDFFRBN $T=722300 366360 0 180 $X=710520 $Y=360940
X692 2693 480 2675 2 1 2670 QDFFRBN $T=724160 305880 0 180 $X=712380 $Y=300460
X693 2676 480 2675 2 1 2669 QDFFRBN $T=724780 285720 0 180 $X=713000 $Y=280300
X694 2696 480 2675 2 1 2620 QDFFRBN $T=727260 295800 1 180 $X=715480 $Y=295420
X695 2700 480 522 2 1 2715 QDFFRBN $T=719200 346200 0 0 $X=719200 $Y=345820
X696 2711 480 2678 2 1 2639 QDFFRBN $T=732840 315960 0 180 $X=721060 $Y=310540
X697 2708 480 520 2 1 2740 QDFFRBN $T=722300 356280 0 0 $X=722300 $Y=355900
X698 2699 480 526 2 1 2704 QDFFRBN $T=722920 265560 0 0 $X=722920 $Y=265180
X699 2718 480 2735 2 1 2729 QDFFRBN $T=725400 336120 0 0 $X=725400 $Y=335740
X700 529 480 522 2 1 510 QDFFRBN $T=737180 366360 0 180 $X=725400 $Y=360940
X701 2721 480 2735 2 1 2755 QDFFRBN $T=726020 346200 1 0 $X=726020 $Y=340780
X702 2722 480 2735 2 1 2746 QDFFRBN $T=726640 305880 1 0 $X=726640 $Y=300460
X703 2723 480 2602 2 1 2751 QDFFRBN $T=727880 285720 1 0 $X=727880 $Y=280300
X704 2725 480 2735 2 1 2757 QDFFRBN $T=729120 305880 0 0 $X=729120 $Y=305500
X705 2783 480 2735 2 1 2716 QDFFRBN $T=747100 336120 0 180 $X=735320 $Y=330700
X706 2759 480 2767 2 1 2795 QDFFRBN $T=740900 305880 1 0 $X=740900 $Y=300460
X707 540 480 2793 2 1 546 QDFFRBN $T=743380 366360 1 0 $X=743380 $Y=360940
X708 2769 480 2767 2 1 2805 QDFFRBN $T=744620 305880 0 0 $X=744620 $Y=305500
X709 2778 480 2793 2 1 553 QDFFRBN $T=747100 356280 0 0 $X=747100 $Y=355900
X710 2785 480 2810 2 1 2798 QDFFRBN $T=748960 326040 0 0 $X=748960 $Y=325660
X711 2787 480 2810 2 1 2821 QDFFRBN $T=749580 356280 1 0 $X=749580 $Y=350860
X712 2808 557 2833 2 1 2844 QDFFRBN $T=757640 295800 0 0 $X=757640 $Y=295420
X713 2811 557 2810 2 1 2776 QDFFRBN $T=757640 326040 1 0 $X=757640 $Y=320620
X714 2814 557 2767 2 1 2845 QDFFRBN $T=758260 305880 1 0 $X=758260 $Y=300460
X715 2824 557 2810 2 1 2834 QDFFRBN $T=763840 326040 0 0 $X=763840 $Y=325660
X716 2832 557 2793 2 1 2860 QDFFRBN $T=765080 356280 1 0 $X=765080 $Y=350860
X717 2861 557 2793 2 1 564 QDFFRBN $T=778100 356280 1 180 $X=766320 $Y=355900
X718 2851 557 2833 2 1 2885 QDFFRBN $T=771900 295800 0 0 $X=771900 $Y=295420
X719 2853 557 2833 2 1 2874 QDFFRBN $T=772520 305880 1 0 $X=772520 $Y=300460
X720 2876 557 2793 2 1 575 QDFFRBN $T=791120 356280 0 180 $X=779340 $Y=350860
X721 2871 557 2909 2 1 2914 QDFFRBN $T=784300 315960 0 0 $X=784300 $Y=315580
X722 2891 557 2833 2 1 2924 QDFFRBN $T=785540 305880 1 0 $X=785540 $Y=300460
X723 2892 557 2909 2 1 2897 QDFFRBN $T=785540 315960 1 0 $X=785540 $Y=310540
X724 2899 557 2915 2 1 2925 QDFFRBN $T=788020 326040 1 0 $X=788020 $Y=320620
X725 2900 557 2915 2 1 2928 QDFFRBN $T=789260 336120 1 0 $X=789260 $Y=330700
X726 2939 557 582 2 1 2910 QDFFRBN $T=805380 346200 1 180 $X=793600 $Y=345820
X727 2920 557 582 2 1 2896 QDFFRBN $T=805380 356280 0 180 $X=793600 $Y=350860
X728 2952 557 2833 2 1 2926 QDFFRBN $T=811580 295800 1 180 $X=799800 $Y=295420
X729 2936 557 2915 2 1 2886 QDFFRBN $T=802280 346200 1 0 $X=802280 $Y=340780
X730 2932 557 2909 2 1 2940 QDFFRBN $T=802900 326040 1 0 $X=802900 $Y=320620
X731 2938 557 2909 2 1 2951 QDFFRBN $T=803520 315960 1 0 $X=803520 $Y=310540
X732 2934 557 2833 2 1 2962 QDFFRBN $T=805380 295800 1 0 $X=805380 $Y=290380
X733 2953 557 582 2 1 600 QDFFRBN $T=819640 356280 0 180 $X=807860 $Y=350860
X734 2949 557 2915 2 1 2961 QDFFRBN $T=808480 346200 0 0 $X=808480 $Y=345820
X735 620 557 633 2 1 640 QDFFRBN $T=812200 366360 1 0 $X=812200 $Y=360940
X736 2966 557 2993 2 1 2973 QDFFRBN $T=821500 326040 1 0 $X=821500 $Y=320620
X737 635 557 633 2 1 639 QDFFRBN $T=822120 356280 1 0 $X=822120 $Y=350860
X738 2979 557 2915 2 1 3005 QDFFRBN $T=823360 346200 0 0 $X=823360 $Y=345820
X739 661 557 633 2 1 644 QDFFRBN $T=837000 366360 0 180 $X=825220 $Y=360940
X740 2983 659 2909 2 1 2977 QDFFRBN $T=837620 315960 1 180 $X=825840 $Y=315580
X741 3007 659 2909 2 1 2985 QDFFRBN $T=842580 305880 1 180 $X=830800 $Y=305500
X742 663 557 633 2 1 680 QDFFRBN $T=837000 356280 0 0 $X=837000 $Y=355900
X743 665 557 633 2 1 688 QDFFRBN $T=837620 366360 1 0 $X=837620 $Y=360940
X744 3013 669 679 2 1 3023 QDFFRBN $T=838240 346200 0 0 $X=838240 $Y=345820
X745 3009 669 2915 2 1 3003 QDFFRBN $T=839480 346200 1 0 $X=839480 $Y=340780
X746 3036 669 2993 2 1 2942 QDFFRBN $T=856220 326040 0 180 $X=844440 $Y=320620
X747 3035 659 3024 2 1 3018 QDFFRBN $T=856840 305880 1 180 $X=845060 $Y=305500
X748 3022 659 3024 2 1 2997 QDFFRBN $T=858080 315960 0 180 $X=846300 $Y=310540
X749 702 669 679 2 1 683 QDFFRBN $T=861180 356280 1 180 $X=849400 $Y=355900
X750 3030 669 2993 2 1 3056 QDFFRBN $T=850640 326040 0 0 $X=850640 $Y=325660
X751 3062 669 2993 2 1 3037 QDFFRBN $T=866140 336120 0 180 $X=854360 $Y=330700
X752 3058 669 679 2 1 3039 QDFFRBN $T=866760 346200 0 180 $X=854980 $Y=340780
X753 3053 659 3024 2 1 3042 QDFFRBN $T=860560 305880 0 0 $X=860560 $Y=305500
X754 3027 659 3024 2 1 3081 QDFFRBN $T=860560 315960 0 0 $X=860560 $Y=315580
X755 3080 659 3061 2 1 3043 QDFFRBN $T=872960 295800 0 180 $X=861180 $Y=290380
X756 3091 669 679 2 1 671 QDFFRBN $T=874820 356280 1 180 $X=863040 $Y=355900
X757 715 669 679 2 1 699 QDFFRBN $T=875440 366360 0 180 $X=863660 $Y=360940
X758 3057 659 3061 2 1 3038 QDFFRBN $T=864280 285720 0 0 $X=864280 $Y=285340
X759 3051 669 679 2 1 3040 QDFFRBN $T=877300 356280 0 180 $X=865520 $Y=350860
X760 3064 659 3090 2 1 3071 QDFFRBN $T=866760 305880 1 0 $X=866760 $Y=300460
X761 3075 669 3085 2 1 3077 QDFFRBN $T=869240 336120 0 0 $X=869240 $Y=335740
X762 3076 669 3085 2 1 3092 QDFFRBN $T=869240 346200 1 0 $X=869240 $Y=340780
X763 3109 659 3061 2 1 2779 QDFFRBN $T=882880 275640 1 180 $X=871100 $Y=275260
X764 3113 659 3090 2 1 3102 QDFFRBN $T=892180 305880 0 180 $X=880400 $Y=300460
X765 3097 659 3090 2 1 609 QDFFRBN $T=892180 315960 0 180 $X=880400 $Y=310540
X766 3126 659 3090 2 1 2903 QDFFRBN $T=892800 305880 1 180 $X=881020 $Y=305500
X767 3124 659 3061 2 1 3002 QDFFRBN $T=894040 295800 0 180 $X=882260 $Y=290380
X768 3130 669 3119 2 1 3089 QDFFRBN $T=894660 326040 0 180 $X=882880 $Y=320620
X769 3131 669 3119 2 1 3083 QDFFRBN $T=894660 326040 1 180 $X=882880 $Y=325660
X770 3122 669 3119 2 1 3096 QDFFRBN $T=895280 336120 1 180 $X=883500 $Y=335740
X771 3114 669 3125 2 1 3133 QDFFRBN $T=883500 346200 1 0 $X=883500 $Y=340780
X772 3098 659 3061 2 1 3107 QDFFRBN $T=884120 285720 1 0 $X=884120 $Y=280300
X773 3115 669 732 2 1 3108 QDFFRBN $T=897140 356280 1 180 $X=885360 $Y=355900
X774 3146 659 3129 2 1 593 QDFFRBN $T=901480 315960 1 180 $X=889700 $Y=315580
X775 3127 669 738 2 1 3112 QDFFRBN $T=891560 356280 1 0 $X=891560 $Y=350860
X776 3151 659 3129 2 1 606 QDFFRBN $T=905200 305880 0 180 $X=893420 $Y=300460
X777 3143 659 3137 2 1 2719 QDFFRBN $T=905820 275640 0 180 $X=894040 $Y=270220
X778 3123 659 3129 2 1 2963 QDFFRBN $T=905820 295800 1 180 $X=894040 $Y=295420
X779 3153 659 3137 2 1 3128 QDFFRBN $T=906440 275640 1 180 $X=894660 $Y=275260
X780 3101 659 3061 2 1 2989 QDFFRBN $T=907680 285720 1 180 $X=895900 $Y=285340
X781 3162 669 3125 2 1 3139 QDFFRBN $T=909540 336120 1 180 $X=897760 $Y=335740
X782 3141 659 3129 2 1 3176 QDFFRBN $T=898380 315960 1 0 $X=898380 $Y=310540
X783 3163 669 3125 2 1 3140 QDFFRBN $T=910160 346200 0 180 $X=898380 $Y=340780
X784 3142 659 3129 2 1 3173 QDFFRBN $T=899000 305880 0 0 $X=899000 $Y=305500
X785 3166 659 744 2 1 720 QDFFRBN $T=913260 265560 0 180 $X=901480 $Y=260140
X786 3170 669 738 2 1 746 QDFFRBN $T=916360 356280 0 180 $X=904580 $Y=350860
X787 3161 659 3137 2 1 3186 QDFFRBN $T=907680 285720 1 0 $X=907680 $Y=280300
X788 3168 659 3137 2 1 3199 QDFFRBN $T=909540 285720 0 0 $X=909540 $Y=285340
X789 3169 669 759 2 1 3184 QDFFRBN $T=909540 356280 0 0 $X=909540 $Y=355900
X790 751 669 759 2 1 765 QDFFRBN $T=911400 366360 1 0 $X=911400 $Y=360940
X791 3179 669 3125 2 1 3134 QDFFRBN $T=912020 336120 1 0 $X=912020 $Y=330700
X792 3198 669 3125 2 1 753 QDFFRBN $T=923800 346200 0 180 $X=912020 $Y=340780
X793 3182 659 766 2 1 3172 QDFFRBN $T=915120 265560 0 0 $X=915120 $Y=265180
X794 3216 659 3197 2 1 3189 QDFFRBN $T=930000 315960 0 180 $X=918220 $Y=310540
X795 3192 659 3209 2 1 774 QDFFRBN $T=920080 275640 1 0 $X=920080 $Y=270220
X796 3202 659 3209 2 1 3233 QDFFRBN $T=923800 285720 0 0 $X=923800 $Y=285340
X797 3207 659 3209 2 1 3235 QDFFRBN $T=925040 295800 0 0 $X=925040 $Y=295420
X798 3211 659 3221 2 1 3240 QDFFRBN $T=926280 326040 1 0 $X=926280 $Y=320620
X799 3217 669 3221 2 1 3188 QDFFRBN $T=938060 336120 1 180 $X=926280 $Y=335740
X800 3213 659 3236 2 1 3243 QDFFRBN $T=927520 285720 1 0 $X=927520 $Y=280300
X801 3214 669 3234 2 1 768 QDFFRBN $T=927520 346200 0 0 $X=927520 $Y=345820
X802 3225 659 3221 2 1 3227 QDFFRBN $T=931240 315960 0 0 $X=931240 $Y=315580
X803 3228 669 759 2 1 796 QDFFRBN $T=932480 356280 0 0 $X=932480 $Y=355900
X804 3226 659 3209 2 1 3229 QDFFRBN $T=934960 275640 1 0 $X=934960 $Y=270220
X805 3252 801 3234 2 1 787 QDFFRBN $T=949220 346200 0 180 $X=937440 $Y=340780
X806 3241 659 766 2 1 803 QDFFRBN $T=938060 265560 1 0 $X=938060 $Y=260140
X807 3261 659 3236 2 1 3239 QDFFRBN $T=951700 305880 0 180 $X=939920 $Y=300460
X808 3244 659 3221 2 1 3264 QDFFRBN $T=939920 315960 1 0 $X=939920 $Y=310540
X809 3231 801 3234 2 1 750 QDFFRBN $T=951700 336120 1 180 $X=939920 $Y=335740
X810 808 801 795 2 1 793 QDFFRBN $T=951700 366360 0 180 $X=939920 $Y=360940
X811 3245 659 3236 2 1 3255 QDFFRBN $T=941780 285720 1 0 $X=941780 $Y=280300
X812 3247 659 3236 2 1 3266 QDFFRBN $T=942400 295800 1 0 $X=942400 $Y=290380
X813 3304 801 3277 2 1 3248 QDFFRBN $T=965340 315960 1 180 $X=953560 $Y=315580
X814 3260 659 3221 2 1 3281 QDFFRBN $T=953560 326040 1 0 $X=953560 $Y=320620
X815 3287 801 3234 2 1 3259 QDFFRBN $T=965340 346200 0 180 $X=953560 $Y=340780
X816 3292 801 822 2 1 814 QDFFRBN $T=965340 366360 0 180 $X=953560 $Y=360940
X817 3296 801 3277 2 1 3262 QDFFRBN $T=966580 326040 1 180 $X=954800 $Y=325660
X818 3280 801 3234 2 1 3272 QDFFRBN $T=966580 336120 1 180 $X=954800 $Y=335740
X819 3290 801 822 2 1 3273 QDFFRBN $T=966580 356280 0 180 $X=954800 $Y=350860
X820 3320 801 822 2 1 3269 QDFFRBN $T=978360 356280 0 180 $X=966580 $Y=350860
X821 3332 801 3277 2 1 3249 QDFFRBN $T=980220 336120 1 180 $X=968440 $Y=335740
X822 3348 801 3221 2 1 3250 QDFFRBN $T=980840 326040 1 180 $X=969060 $Y=325660
X823 3339 801 3277 2 1 3263 QDFFRBN $T=981460 336120 0 180 $X=969680 $Y=330700
X824 3333 801 869 2 1 3365 QDFFRBN $T=978360 346200 1 0 $X=978360 $Y=340780
X825 3334 801 869 2 1 3349 QDFFRBN $T=978360 356280 1 0 $X=978360 $Y=350860
X826 3415 801 869 2 1 3383 QDFFRBN $T=1005020 346200 0 180 $X=993240 $Y=340780
X827 3388 801 869 2 1 3362 QDFFRBN $T=994480 356280 0 0 $X=994480 $Y=355900
X828 3433 801 3432 2 1 3421 QDFFRBN $T=1008740 346200 1 0 $X=1008740 $Y=340780
X829 3463 801 3432 2 1 3441 QDFFRBN $T=1021140 336120 1 180 $X=1009360 $Y=335740
X830 3481 659 915 2 1 910 QDFFRBN $T=1026100 265560 0 180 $X=1014320 $Y=260140
X831 922 659 915 2 1 3420 QDFFRBN $T=1026720 275640 0 180 $X=1014940 $Y=270220
X832 928 659 915 2 1 3409 QDFFRBN $T=1027960 275640 1 180 $X=1016180 $Y=275260
X833 3470 801 3485 2 1 3475 QDFFRBN $T=1018660 356280 0 0 $X=1018660 $Y=355900
X834 3472 801 3485 2 1 947 QDFFRBN $T=1024240 346200 0 0 $X=1024240 $Y=345820
X835 954 905 915 2 1 3411 QDFFRBN $T=1041600 275640 1 180 $X=1029820 $Y=275260
X836 3520 905 3485 2 1 3491 QDFFRBN $T=1041600 346200 0 180 $X=1029820 $Y=340780
X837 956 953 943 2 1 937 QDFFRBN $T=1042220 356280 1 180 $X=1030440 $Y=355900
X838 3505 905 3486 2 1 3482 QDFFRBN $T=1031680 295800 0 0 $X=1031680 $Y=295420
X839 3532 905 3486 2 1 3359 QDFFRBN $T=1044700 285720 0 180 $X=1032920 $Y=280300
X840 3502 905 3529 2 1 3540 QDFFRBN $T=1032920 305880 1 0 $X=1032920 $Y=300460
X841 3517 905 3530 2 1 3537 QDFFRBN $T=1034780 295800 1 0 $X=1034780 $Y=290380
X842 3546 905 3485 2 1 952 QDFFRBN $T=1050280 356280 0 180 $X=1038500 $Y=350860
X843 3533 905 3551 2 1 3560 QDFFRBN $T=1042840 326040 1 0 $X=1042840 $Y=320620
X844 3534 905 3554 2 1 979 QDFFRBN $T=1044080 346200 1 0 $X=1044080 $Y=340780
X845 3536 905 3551 2 1 3563 QDFFRBN $T=1044700 336120 1 0 $X=1044700 $Y=330700
X846 968 953 943 2 1 988 QDFFRBN $T=1044700 356280 0 0 $X=1044700 $Y=355900
X847 3538 905 3530 2 1 3567 QDFFRBN $T=1045940 305880 0 0 $X=1045940 $Y=305500
X848 3544 905 3530 2 1 3576 QDFFRBN $T=1047800 305880 1 0 $X=1047800 $Y=300460
X849 3594 905 3529 2 1 3548 QDFFRBN $T=1062060 285720 0 180 $X=1050280 $Y=280300
X850 3587 905 3530 2 1 3531 QDFFRBN $T=1062060 295800 0 180 $X=1050280 $Y=290380
X851 3586 905 3554 2 1 3557 QDFFRBN $T=1066400 346200 1 180 $X=1054620 $Y=345820
X852 3564 905 3529 2 1 3581 QDFFRBN $T=1055860 275640 0 0 $X=1055860 $Y=275260
X853 3572 905 3554 2 1 3612 QDFFRBN $T=1057720 336120 0 0 $X=1057720 $Y=335740
X854 3591 905 943 2 1 3561 QDFFRBN $T=1075080 356280 0 180 $X=1063300 $Y=350860
X855 1005 905 943 2 1 996 QDFFRBN $T=1076320 366360 0 180 $X=1064540 $Y=360940
X856 3648 905 3554 2 1 3606 QDFFRBN $T=1079420 346200 0 180 $X=1067640 $Y=340780
X857 3653 905 3529 2 1 3611 QDFFRBN $T=1080660 265560 1 180 $X=1068880 $Y=265180
X858 3664 905 3551 2 1 3617 QDFFRBN $T=1083760 336120 1 180 $X=1071980 $Y=335740
X859 3685 905 3554 2 1 3665 QDFFRBN $T=1092440 346200 1 180 $X=1080660 $Y=345820
X860 3668 905 3551 2 1 3667 QDFFRBN $T=1081280 336120 1 0 $X=1081280 $Y=330700
X861 3673 905 3529 2 1 3682 QDFFRBN $T=1083140 265560 0 0 $X=1083140 $Y=265180
X862 3702 905 3554 2 1 3671 QDFFRBN $T=1094920 346200 0 180 $X=1083140 $Y=340780
X863 3701 905 3692 2 1 3683 QDFFRBN $T=1098640 285720 1 180 $X=1086860 $Y=285340
X864 3722 905 3692 2 1 3605 QDFFRBN $T=1099880 295800 0 180 $X=1088100 $Y=290380
X865 3688 905 3715 2 1 3626 QDFFRBN $T=1088100 305880 0 0 $X=1088100 $Y=305500
X866 3675 905 3551 2 1 3652 QDFFRBN $T=1101120 315960 1 180 $X=1089340 $Y=315580
X867 3712 905 3715 2 1 3743 QDFFRBN $T=1094920 305880 1 0 $X=1094920 $Y=300460
X868 3713 905 3737 2 1 3718 QDFFRBN $T=1094920 336120 1 0 $X=1094920 $Y=330700
X869 3742 905 3721 2 1 3693 QDFFRBN $T=1106700 356280 1 180 $X=1094920 $Y=355900
X870 3728 905 3721 2 1 3660 QDFFRBN $T=1107320 346200 1 180 $X=1095540 $Y=345820
X871 3745 905 3692 2 1 3731 QDFFRBN $T=1112900 285720 1 180 $X=1101120 $Y=285340
X872 3717 905 3721 2 1 3694 QDFFRBN $T=1113520 356280 0 180 $X=1101740 $Y=350860
X873 3740 905 1038 2 1 3771 QDFFRBN $T=1103600 265560 0 0 $X=1103600 $Y=265180
X874 3760 905 3721 2 1 3744 QDFFRBN $T=1116000 346200 0 180 $X=1104220 $Y=340780
X875 3800 905 1038 2 1 3754 QDFFRBN $T=1127780 275640 1 180 $X=1116000 $Y=275260
X876 3789 905 3715 2 1 3779 QDFFRBN $T=1116000 285720 0 0 $X=1116000 $Y=285340
X877 3793 905 3737 2 1 3756 QDFFRBN $T=1127780 315960 0 180 $X=1116000 $Y=310540
X878 3790 905 1038 2 1 3801 QDFFRBN $T=1116620 275640 1 0 $X=1116620 $Y=270220
X879 3782 905 3715 2 1 3776 QDFFRBN $T=1128400 305880 0 180 $X=1116620 $Y=300460
X880 3727 905 3737 2 1 3802 QDFFRBN $T=1116620 315960 0 0 $X=1116620 $Y=315580
X881 3791 905 3737 2 1 3748 QDFFRBN $T=1116620 326040 1 0 $X=1116620 $Y=320620
X882 3786 905 3737 2 1 3741 QDFFRBN $T=1116620 336120 0 0 $X=1116620 $Y=335740
X883 3778 905 3721 2 1 3764 QDFFRBN $T=1128400 356280 0 180 $X=1116620 $Y=350860
X884 3794 905 1046 2 1 3768 QDFFRBN $T=1128400 366360 0 180 $X=1116620 $Y=360940
X885 2716 1 2 2728 2729 2707 1070 ICV_4 $T=725400 336120 1 0 $X=725400 $Y=330700
X886 2896 1 2 2912 599 605 1070 ICV_4 $T=794840 356280 0 0 $X=794840 $Y=355900
X887 600 1 2 2943 612 622 1070 ICV_4 $T=803520 336120 1 0 $X=803520 $Y=330700
X888 610 1 2 615 616 625 1070 ICV_4 $T=806000 356280 0 0 $X=806000 $Y=355900
X889 623 1 2 628 630 636 1070 ICV_4 $T=813440 336120 1 0 $X=813440 $Y=330700
X890 671 1 2 3021 3023 3029 1070 ICV_4 $T=841340 356280 1 0 $X=841340 $Y=350860
X891 687 1 2 693 3042 3050 1070 ICV_4 $T=850640 305880 1 0 $X=850640 $Y=300460
X892 688 1 2 694 683 704 1070 ICV_4 $T=851260 366360 1 0 $X=851260 $Y=360940
X893 3040 1 2 3048 3039 3049 1070 ICV_4 $T=854980 336120 0 0 $X=854980 $Y=335740
X894 699 1 2 707 3037 3067 1070 ICV_4 $T=858080 315960 1 0 $X=858080 $Y=310540
X895 3071 1 2 3070 3078 3075 1070 ICV_4 $T=868000 315960 1 0 $X=868000 $Y=310540
X896 716 1 2 725 3108 3103 1070 ICV_4 $T=876060 366360 1 0 $X=876060 $Y=360940
X897 3096 1 2 3117 3112 3116 1070 ICV_4 $T=885360 336120 1 0 $X=885360 $Y=330700
X898 3188 1 2 3201 780 785 1070 ICV_4 $T=925660 326040 0 0 $X=925660 $Y=325660
X899 772 1 2 3212 782 788 1070 ICV_4 $T=927520 356280 1 0 $X=927520 $Y=350860
X900 821 1 2 828 830 836 1070 ICV_4 $T=956660 356280 0 0 $X=956660 $Y=355900
X901 3540 1 2 3484 3556 3538 1070 ICV_4 $T=1049040 295800 0 0 $X=1049040 $Y=295420
X902 1010 1 2 1016 3665 3676 1070 ICV_4 $T=1078800 356280 0 0 $X=1078800 $Y=355900
X903 3671 1 2 3687 1023 1026 1070 ICV_4 $T=1088100 336120 0 0 $X=1088100 $Y=335740
X904 1028 1 2 1031 3694 3703 1070 ICV_4 $T=1100500 336120 0 0 $X=1100500 $Y=335740
X905 3764 1 2 3757 1051 1054 1070 ICV_4 $T=1118480 356280 0 0 $X=1118480 $Y=355900
X906 1372 100 2 1 1414 1406 MUX2 $T=318680 366360 1 0 $X=318680 $Y=360940
X907 1389 100 2 1 1438 1431 MUX2 $T=323020 346200 1 0 $X=323020 $Y=340780
X908 1400 100 2 1 1385 1432 MUX2 $T=324880 356280 1 0 $X=324880 $Y=350860
X909 1410 1435 2 1 1454 1455 MUX2 $T=329840 336120 0 0 $X=329840 $Y=335740
X910 1450 1435 2 1 1466 1461 MUX2 $T=332320 315960 0 0 $X=332320 $Y=315580
X911 1445 1435 2 1 1468 1472 MUX2 $T=332940 305880 0 0 $X=332940 $Y=305500
X912 1467 1435 2 1 1465 1460 MUX2 $T=336660 295800 0 0 $X=336660 $Y=295420
X913 1458 108 2 1 1495 1483 MUX2 $T=337900 275640 1 0 $X=337900 $Y=270220
X914 1479 1435 2 1 1493 1492 MUX2 $T=340380 295800 1 0 $X=340380 $Y=290380
X915 1471 108 2 1 1510 1509 MUX2 $T=346580 285720 1 0 $X=346580 $Y=280300
X916 2174 341 2 1 323 345 MUX2 $T=554280 366360 1 0 $X=554280 $Y=360940
X917 2681 2677 2 1 2643 2671 MUX2 $T=714860 326040 0 0 $X=714860 $Y=325660
X918 556 554 2 1 2778 548 MUX2 $T=759500 366360 0 180 $X=755160 $Y=360940
X919 570 569 2 1 2861 573 MUX2 $T=773760 366360 1 0 $X=773760 $Y=360940
X920 2868 554 2 1 2876 573 MUX2 $T=778100 366360 1 0 $X=778100 $Y=360940
X921 2887 554 2 1 580 579 MUX2 $T=786780 366360 0 180 $X=782440 $Y=360940
X922 2912 569 2 1 2920 579 MUX2 $T=794220 366360 1 0 $X=794220 $Y=360940
X923 2924 2935 2 1 596 2874 MUX2 $T=802280 305880 1 180 $X=797940 $Y=305500
X924 2933 554 2 1 2939 608 MUX2 $T=802280 366360 1 0 $X=802280 $Y=360940
X925 2943 569 2 1 2953 608 MUX2 $T=806620 366360 1 0 $X=806620 $Y=360940
X926 2962 2935 2 1 619 2897 MUX2 $T=817780 295800 1 180 $X=813440 $Y=295420
X927 2885 2964 2 1 624 2940 MUX2 $T=820260 305880 1 180 $X=815920 $Y=305500
X928 3029 3044 2 1 3013 690 MUX2 $T=855600 356280 0 180 $X=851260 $Y=350860
X929 3049 3044 2 1 3058 708 MUX2 $T=859940 346200 0 0 $X=859940 $Y=345820
X930 3048 710 2 1 3051 690 MUX2 $T=864280 356280 0 180 $X=859940 $Y=350860
X931 3067 710 2 1 3062 708 MUX2 $T=868620 346200 1 180 $X=864280 $Y=345820
X932 3094 710 2 1 3076 714 MUX2 $T=876680 346200 1 180 $X=872340 $Y=345820
X933 3102 2982 2 1 718 3038 MUX2 $T=880400 295800 0 180 $X=876060 $Y=290380
X934 3021 724 2 1 3091 714 MUX2 $T=880400 356280 1 180 $X=876060 $Y=355900
X935 3103 726 2 1 3115 730 MUX2 $T=880400 356280 1 0 $X=880400 $Y=350860
X936 3107 2982 2 1 3082 2719 MUX2 $T=887220 275640 1 180 $X=882880 $Y=275260
X937 3116 710 2 1 3127 730 MUX2 $T=884740 356280 1 0 $X=884740 $Y=350860
X938 3117 3044 2 1 3122 714 MUX2 $T=885360 346200 0 0 $X=885360 $Y=345820
X939 3128 2982 2 1 717 2779 MUX2 $T=892800 275640 1 180 $X=888460 $Y=275260
X940 3132 3044 2 1 3114 737 MUX2 $T=893420 346200 0 0 $X=893420 $Y=345820
X941 3150 724 2 1 3170 737 MUX2 $T=903960 366360 1 0 $X=903960 $Y=360940
X942 3156 3145 2 1 3163 737 MUX2 $T=906440 346200 0 0 $X=906440 $Y=345820
X943 3185 3145 2 1 3169 754 MUX2 $T=917600 346200 1 180 $X=913260 $Y=345820
X944 3187 758 2 1 3198 754 MUX2 $T=917600 346200 0 0 $X=917600 $Y=345820
X945 3201 726 2 1 3217 754 MUX2 $T=923800 346200 1 0 $X=923800 $Y=340780
X946 3319 3291 2 1 854 853 MUX2 $T=974020 366360 1 0 $X=974020 $Y=360940
X947 3562 3549 2 1 3534 984 MUX2 $T=1058340 356280 0 180 $X=1054000 $Y=350860
X948 3574 992 2 1 3586 984 MUX2 $T=1058340 356280 1 0 $X=1058340 $Y=350860
X949 3575 951 2 1 3591 984 MUX2 $T=1058960 356280 0 0 $X=1058960 $Y=355900
X950 3640 1004 2 1 3648 1012 MUX2 $T=1075080 356280 1 0 $X=1075080 $Y=350860
X951 3676 1004 2 1 3685 1020 MUX2 $T=1083760 356280 1 0 $X=1083760 $Y=350860
X952 3687 3549 2 1 3702 1020 MUX2 $T=1088100 356280 1 0 $X=1088100 $Y=350860
X953 3704 3549 2 1 3728 1012 MUX2 $T=1093060 356280 1 0 $X=1093060 $Y=350860
X954 3703 3549 2 1 3717 1025 MUX2 $T=1093060 366360 1 0 $X=1093060 $Y=360940
X955 3709 1004 2 1 3742 1025 MUX2 $T=1098020 366360 1 0 $X=1098020 $Y=360940
X956 3757 951 2 1 3778 1012 MUX2 $T=1109180 356280 0 0 $X=1109180 $Y=355900
X957 3780 992 2 1 3794 1012 MUX2 $T=1114140 356280 0 0 $X=1114140 $Y=355900
X958 2012 1976 2005 1989 1 1954 2 AOI22S $T=510880 356280 0 180 $X=507160 $Y=350860
X959 2012 1990 2007 1989 1 1976 2 AOI22S $T=514600 346200 1 180 $X=510880 $Y=345820
X960 2012 2023 2035 293 1 1990 2 AOI22S $T=518320 346200 1 180 $X=514600 $Y=345820
X961 2004 2025 2031 2023 1 293 2 AOI22S $T=519560 346200 0 180 $X=515840 $Y=340780
X962 2012 2047 2051 1989 1 2023 2 AOI22S $T=525140 356280 0 180 $X=521420 $Y=350860
X963 2043 2034 299 301 1 305 2 AOI22S $T=521420 366360 1 0 $X=521420 $Y=360940
X964 2004 1989 2049 2023 1 2012 2 AOI22S $T=523280 346200 1 0 $X=523280 $Y=340780
X965 303 304 2052 301 1 305 2 AOI22S $T=524520 356280 0 0 $X=524520 $Y=355900
X966 2012 2061 2065 1989 1 2047 2 AOI22S $T=529480 356280 0 180 $X=525760 $Y=350860
X967 2067 307 308 301 1 305 2 AOI22S $T=529480 366360 0 180 $X=525760 $Y=360940
X968 288 311 2078 301 1 305 2 AOI22S $T=532580 356280 1 180 $X=528860 $Y=355900
X969 2061 2084 2079 2074 1 2089 2 AOI22S $T=531340 336120 1 0 $X=531340 $Y=330700
X970 2089 2090 2098 2074 1 2084 2 AOI22S $T=535060 336120 0 0 $X=535060 $Y=335740
X971 2090 2111 2121 2074 1 2089 2 AOI22S $T=542500 336120 1 180 $X=538780 $Y=335740
X972 2089 2137 2142 2074 1 2111 2 AOI22S $T=545600 336120 0 0 $X=545600 $Y=335740
X973 2162 2149 2165 2169 1 2137 2 AOI22S $T=549320 346200 1 0 $X=549320 $Y=340780
X974 2089 2177 2176 2074 1 2168 2 AOI22S $T=553660 336120 0 0 $X=553660 $Y=335740
X975 2149 2168 2181 2169 1 2162 2 AOI22S $T=554280 336120 1 0 $X=554280 $Y=330700
X976 2177 2190 2189 2169 1 2162 2 AOI22S $T=558000 336120 1 0 $X=558000 $Y=330700
X977 2225 350 2217 2180 1 2162 2 AOI22S $T=564820 336120 1 180 $X=561100 $Y=335740
X978 2212 2133 2193 350 1 2216 2 AOI22S $T=562960 356280 1 0 $X=562960 $Y=350860
X979 2218 2133 2207 358 1 2216 2 AOI22S $T=563580 356280 0 0 $X=563580 $Y=355900
X980 350 363 2204 365 1 367 2 AOI22S $T=566680 366360 1 0 $X=566680 $Y=360940
X981 2218 363 2203 358 1 367 2 AOI22S $T=567300 356280 0 0 $X=567300 $Y=355900
X982 2216 2225 2227 367 1 2242 2 AOI22S $T=567920 346200 1 0 $X=567920 $Y=340780
X983 2216 2242 2226 2200 1 2190 2 AOI22S $T=570400 336120 0 0 $X=570400 $Y=335740
X984 2242 2201 2248 2216 1 367 2 AOI22S $T=571640 346200 1 0 $X=571640 $Y=340780
X985 2169 2218 2235 2200 1 2212 2 AOI22S $T=575360 336120 1 0 $X=575360 $Y=330700
X986 558 585 587 2896 1 578 2 AOI22S $T=790500 366360 0 180 $X=786780 $Y=360940
X987 558 585 597 600 1 2910 2 AOI22S $T=798560 366360 1 0 $X=798560 $Y=360940
X988 2982 2844 638 2964 1 2973 2 AOI22S $T=824600 305880 1 180 $X=820880 $Y=305500
X989 2982 2985 649 2964 1 2977 2 AOI22S $T=828320 305880 1 180 $X=824600 $Y=305500
X990 700 3041 696 3039 1 3037 2 AOI22S $T=857460 346200 1 180 $X=853740 $Y=345820
X991 700 3041 697 3023 1 3040 2 AOI22S $T=859320 356280 0 180 $X=855600 $Y=350860
X992 2982 3002 713 3046 1 3071 2 AOI22S $T=871100 295800 0 0 $X=871100 $Y=295420
X993 3100 3041 721 3096 1 3092 2 AOI22S $T=880400 346200 1 180 $X=876680 $Y=345820
X994 700 723 727 3108 1 3112 2 AOI22S $T=881020 356280 0 0 $X=881020 $Y=355900
X995 3100 723 743 3133 1 3140 2 AOI22S $T=902100 346200 0 0 $X=902100 $Y=345820
X996 764 723 760 3188 1 3184 2 AOI22S $T=920700 356280 0 180 $X=916980 $Y=350860
X997 764 771 807 3259 1 3269 2 AOI22S $T=951080 346200 0 0 $X=951080 $Y=345820
X998 764 771 815 3272 1 3273 2 AOI22S $T=952940 356280 0 0 $X=952940 $Y=355900
X999 881 876 3361 3365 1 3349 2 AOI22S $T=992620 366360 0 180 $X=988900 $Y=360940
X1000 881 876 3398 3383 1 3362 2 AOI22S $T=998820 366360 1 0 $X=998820 $Y=360940
X1001 901 902 3395 895 1 3421 2 AOI22S $T=1006880 366360 1 0 $X=1006880 $Y=360940
X1002 901 902 3357 909 1 3441 2 AOI22S $T=1011220 366360 1 0 $X=1011220 $Y=360940
X1003 927 925 930 3475 1 3491 2 AOI22S $T=1026720 366360 1 0 $X=1026720 $Y=360940
X1004 3521 3526 3515 962 1 3506 2 AOI22S $T=1041600 275640 1 0 $X=1041600 $Y=270220
X1005 932 986 3566 3555 1 3553 2 AOI22S $T=1056480 275640 0 180 $X=1052760 $Y=270220
X1006 927 985 982 3557 1 3561 2 AOI22S $T=1052760 366360 1 0 $X=1052760 $Y=360940
X1007 993 939 3601 995 1 965 2 AOI22S $T=1063300 265560 0 180 $X=1059580 $Y=260140
X1008 3624 3632 3608 3638 1 3646 2 AOI22S $T=1073840 285720 0 0 $X=1073840 $Y=285340
X1009 3672 1014 1015 3606 1 3660 2 AOI22S $T=1083140 356280 0 180 $X=1079420 $Y=350860
X1010 3672 1014 1018 3665 1 3671 2 AOI22S $T=1083760 366360 1 0 $X=1083760 $Y=360940
X1011 3672 1014 1021 3693 1 3694 2 AOI22S $T=1088100 366360 1 0 $X=1088100 $Y=360940
X1012 3690 3698 3680 3700 1 3659 2 AOI22S $T=1090580 326040 0 0 $X=1090580 $Y=325660
X1013 1032 985 1035 3768 1 3764 2 AOI22S $T=1107940 366360 1 0 $X=1107940 $Y=360940
X1014 14 2 1 1136 BUF1 $T=233120 326040 1 0 $X=233120 $Y=320620
X1015 13 2 1 1137 BUF1 $T=238080 295800 0 0 $X=238080 $Y=295420
X1016 1101 2 1 1139 BUF1 $T=239940 326040 0 0 $X=239940 $Y=325660
X1017 35 2 1 29 BUF1 $T=243660 356280 0 0 $X=243660 $Y=355900
X1018 1524 2 1 1527 BUF1 $T=354020 295800 1 0 $X=354020 $Y=290380
X1019 1619 2 1 1628 BUF1 $T=385640 326040 0 0 $X=385640 $Y=325660
X1020 157 2 1 1655 BUF1 $T=396800 285720 1 0 $X=396800 $Y=280300
X1021 175 2 1 1637 BUF1 $T=399280 356280 0 180 $X=396800 $Y=350860
X1022 1652 2 1 164 BUF1 $T=404240 336120 0 180 $X=401760 $Y=330700
X1023 1607 2 1 166 BUF1 $T=404240 336120 1 180 $X=401760 $Y=335740
X1024 1697 2 1 182 BUF1 $T=407960 265560 0 180 $X=405480 $Y=260140
X1025 1655 2 1 184 BUF1 $T=405480 336120 0 0 $X=405480 $Y=335740
X1026 176 2 1 1691 BUF1 $T=409820 356280 0 180 $X=407340 $Y=350860
X1027 196 2 1 1722 BUF1 $T=424080 326040 0 180 $X=421600 $Y=320620
X1028 1729 2 1 1723 BUF1 $T=425940 315960 0 180 $X=423460 $Y=310540
X1029 205 2 1 1729 BUF1 $T=429040 346200 1 180 $X=426560 $Y=345820
X1030 219 2 1 1731 BUF1 $T=437720 356280 0 180 $X=435240 $Y=350860
X1031 203 2 1 1766 BUF1 $T=442680 295800 1 180 $X=440200 $Y=295420
X1032 231 2 1 1797 BUF1 $T=444540 315960 1 0 $X=444540 $Y=310540
X1033 231 2 1 221 BUF1 $T=450120 295800 0 0 $X=450120 $Y=295420
X1034 227 2 1 1816 BUF1 $T=451360 295800 1 0 $X=451360 $Y=290380
X1035 1825 2 1 239 BUF1 $T=455080 265560 1 0 $X=455080 $Y=260140
X1036 1829 2 1 1825 BUF1 $T=456320 315960 1 0 $X=456320 $Y=310540
X1037 245 2 1 235 BUF1 $T=464380 265560 0 180 $X=461900 $Y=260140
X1038 245 2 1 1836 BUF1 $T=468100 326040 1 180 $X=465620 $Y=325660
X1039 248 2 1 1829 BUF1 $T=465620 366360 1 0 $X=465620 $Y=360940
X1040 1902 2 1 1862 BUF1 $T=481740 305880 1 180 $X=479260 $Y=305500
X1041 268 2 1 270 BUF1 $T=487320 326040 1 180 $X=484840 $Y=325660
X1042 1926 2 1 1921 BUF1 $T=489180 305880 0 0 $X=489180 $Y=305500
X1043 1957 2 1 1924 BUF1 $T=500340 275640 1 180 $X=497860 $Y=275260
X1044 1964 2 1 2002 BUF1 $T=517700 285720 0 180 $X=515220 $Y=280300
X1045 2016 2 1 2036 BUF1 $T=522040 275640 1 0 $X=522040 $Y=270220
X1046 1999 2 1 2010 BUF1 $T=525140 275640 1 180 $X=522660 $Y=275260
X1047 2166 2 1 2046 BUF1 $T=551800 275640 1 180 $X=549320 $Y=275260
X1048 2160 2 1 2126 BUF1 $T=551800 285720 0 180 $X=549320 $Y=280300
X1049 281 2 1 2205 BUF1 $T=558620 315960 1 0 $X=558620 $Y=310540
X1050 1957 2 1 2222 BUF1 $T=570400 326040 1 0 $X=570400 $Y=320620
X1051 2270 2 1 1964 BUF1 $T=581560 315960 0 180 $X=579080 $Y=310540
X1052 371 2 1 2295 BUF1 $T=586520 356280 0 0 $X=586520 $Y=355900
X1053 402 2 1 2244 BUF1 $T=592720 275640 1 180 $X=590240 $Y=275260
X1054 1999 2 1 2313 BUF1 $T=593340 295800 1 0 $X=593340 $Y=290380
X1055 1999 2 1 401 BUF1 $T=593960 275640 0 0 $X=593960 $Y=275260
X1056 2285 2 1 2305 BUF1 $T=594580 265560 0 0 $X=594580 $Y=265180
X1057 2352 2 1 2166 BUF1 $T=603260 285720 0 180 $X=600780 $Y=280300
X1058 2404 2 1 2454 BUF1 $T=630540 336120 1 0 $X=630540 $Y=330700
X1059 402 2 1 2460 BUF1 $T=633020 285720 0 0 $X=633020 $Y=285340
X1060 420 2 1 2462 BUF1 $T=633020 346200 0 0 $X=633020 $Y=345820
X1061 434 2 1 2426 BUF1 $T=636740 336120 1 180 $X=634260 $Y=335740
X1062 429 2 1 2452 BUF1 $T=634260 366360 1 0 $X=634260 $Y=360940
X1063 435 2 1 2425 BUF1 $T=646660 336120 0 0 $X=646660 $Y=335740
X1064 2381 2 1 2352 BUF1 $T=649140 326040 1 0 $X=649140 $Y=320620
X1065 446 2 1 455 BUF1 $T=656580 315960 1 180 $X=654100 $Y=315580
X1066 450 2 1 454 BUF1 $T=657200 295800 1 0 $X=657200 $Y=290380
X1067 442 2 1 457 BUF1 $T=658440 305880 0 0 $X=658440 $Y=305500
X1068 460 2 1 458 BUF1 $T=660920 326040 0 0 $X=660920 $Y=325660
X1069 2547 2 1 474 BUF1 $T=677660 265560 0 180 $X=675180 $Y=260140
X1070 2731 2 1 2741 BUF1 $T=738420 315960 1 0 $X=738420 $Y=310540
X1071 2872 2 1 2883 BUF1 $T=781820 315960 0 0 $X=781820 $Y=315580
X1072 2884 2 1 2889 BUF1 $T=786780 326040 0 0 $X=786780 $Y=325660
X1073 2694 2 1 2917 BUF1 $T=792360 305880 0 0 $X=792360 $Y=305500
X1074 2964 2 1 2935 BUF1 $T=820260 305880 0 180 $X=817780 $Y=300460
X1075 2917 2 1 2972 BUF1 $T=817780 326040 1 0 $X=817780 $Y=320620
X1076 3046 2 1 2964 BUF1 $T=857460 295800 1 180 $X=854980 $Y=295420
X1077 723 2 1 771 BUF1 $T=923800 356280 1 0 $X=923800 $Y=350860
X1078 925 2 1 985 BUF1 $T=1056480 366360 1 0 $X=1056480 $Y=360940
X1079 1535 1 2 1539 BUF1CK $T=358360 305880 0 0 $X=358360 $Y=305500
X1080 245 1 2 1823 BUF1CK $T=463760 295800 1 0 $X=463760 $Y=290380
X1081 270 1 2 1894 BUF1CK $T=486080 326040 0 180 $X=483600 $Y=320620
X1082 300 1 2 2043 BUF1CK $T=521420 356280 0 0 $X=521420 $Y=355900
X1083 309 1 2 2067 BUF1CK $T=529480 366360 1 0 $X=529480 $Y=360940
X1084 2467 1 2 2453 BUF1CK $T=648520 295800 1 180 $X=646040 $Y=295420
X1085 2620 1 2 2613 BUF1CK $T=696880 295800 0 0 $X=696880 $Y=295420
X1086 2685 1 2 2683 BUF1CK $T=716100 346200 1 0 $X=716100 $Y=340780
X1087 2738 1 2 2733 BUF1CK $T=734080 295800 0 0 $X=734080 $Y=295420
X1088 2818 1 2 2804 BUF1CK $T=758880 356280 0 0 $X=758880 $Y=355900
X1089 589 1 2 585 BUF1CK $T=790500 366360 1 0 $X=790500 $Y=360940
X1090 609 1 2 2984 BUF1CK $T=828320 295800 0 0 $X=828320 $Y=295420
X1091 3063 1 2 3054 BUF1CK $T=874820 326040 1 0 $X=874820 $Y=320620
X1092 700 1 2 3100 BUF1CK $T=880400 346200 0 0 $X=880400 $Y=345820
X1093 3164 1 2 3167 BUF1CK $T=908300 295800 1 0 $X=908300 $Y=290380
X1094 3171 1 2 3177 BUF1CK $T=909540 326040 1 0 $X=909540 $Y=320620
X1095 3215 1 2 3220 BUF1CK $T=927520 315960 0 0 $X=927520 $Y=315580
X1096 3242 1 2 3230 BUF1CK $T=944880 305880 0 0 $X=944880 $Y=305500
X1097 786 1 2 857 BUF1CK $T=983940 366360 1 0 $X=983940 $Y=360940
X1098 3563 1 2 3568 BUF1CK $T=1055240 336120 0 0 $X=1055240 $Y=335740
X1099 3611 1 2 1000 BUF1CK $T=1068880 275640 1 0 $X=1068880 $Y=270220
X1100 3605 1 2 3708 BUF1CK $T=1092440 305880 1 0 $X=1092440 $Y=300460
X1101 3731 1 2 3725 BUF1CK $T=1101120 275640 0 0 $X=1101120 $Y=275260
X1102 3735 1 2 3733 BUF1CK $T=1101740 315960 0 0 $X=1101740 $Y=315580
X1103 3743 1 2 3749 BUF1CK $T=1103600 295800 0 0 $X=1103600 $Y=295420
X1104 927 1 2 1032 BUF1CK $T=1105460 366360 1 0 $X=1105460 $Y=360940
X1105 3781 1 2 3788 BUF1CK $T=1117860 305880 0 0 $X=1117860 $Y=305500
X1106 3796 1 2 3795 BUF1CK $T=1125300 295800 0 0 $X=1125300 $Y=295420
X1107 1745 193 1 2 INV2 $T=426560 295800 0 180 $X=424700 $Y=290380
X1108 1782 1745 1 2 INV2 $T=443920 315960 0 180 $X=442060 $Y=310540
X1109 1888 249 1 2 INV2 $T=473060 265560 1 180 $X=471200 $Y=265180
X1110 1888 256 1 2 INV2 $T=474920 265560 0 0 $X=474920 $Y=265180
X1111 284 1926 1 2 INV2 $T=504680 326040 0 180 $X=502820 $Y=320620
X1112 284 2220 1 2 INV2 $T=563580 326040 0 0 $X=563580 $Y=325660
X1113 364 2206 1 2 INV2 $T=568540 326040 0 0 $X=568540 $Y=325660
X1114 2215 2210 1 2 INV2 $T=569160 305880 1 0 $X=569160 $Y=300460
X1115 2246 1957 1 2 INV2 $T=571020 326040 0 0 $X=571020 $Y=325660
X1116 381 2016 1 2 INV2 $T=581560 326040 1 0 $X=581560 $Y=320620
X1117 381 2285 1 2 INV2 $T=583420 326040 1 0 $X=583420 $Y=320620
X1118 387 2270 1 2 INV2 $T=584660 336120 0 0 $X=584660 $Y=335740
X1119 413 2381 1 2 INV2 $T=610080 336120 0 0 $X=610080 $Y=335740
X1120 445 2198 1 2 INV2 $T=641700 275640 1 180 $X=639840 $Y=275260
X1121 440 2251 1 2 INV2 $T=646040 275640 1 0 $X=646040 $Y=270220
X1122 452 442 1 2 INV2 $T=651620 315960 0 0 $X=651620 $Y=315580
X1123 2548 443 1 2 INV2 $T=665260 285720 0 180 $X=663400 $Y=280300
X1124 462 2548 1 2 INV2 $T=663400 356280 1 0 $X=663400 $Y=350860
X1125 3195 764 1 2 INV2 $T=920700 356280 1 0 $X=920700 $Y=350860
X1126 3661 3672 1 2 INV2 $T=1080660 366360 1 0 $X=1080660 $Y=360940
X1127 197 1715 1 2 BUF2 $T=425320 315960 0 0 $X=425320 $Y=315580
X1128 216 1749 1 2 BUF2 $T=432760 305880 0 0 $X=432760 $Y=305500
X1129 222 1782 1 2 BUF2 $T=439580 366360 1 0 $X=439580 $Y=360940
X1130 1894 1869 1 2 BUF2 $T=478640 326040 0 180 $X=475540 $Y=320620
X1131 1921 278 1 2 BUF2 $T=494140 275640 0 0 $X=494140 $Y=275260
X1132 1957 282 1 2 BUF2 $T=509020 275640 0 180 $X=505920 $Y=270220
X1133 2206 281 1 2 BUF2 $T=561100 315960 1 0 $X=561100 $Y=310540
X1134 2269 1999 1 2 BUF2 $T=581560 315960 1 0 $X=581560 $Y=310540
X1135 2265 2309 1 2 BUF2 $T=587140 336120 0 0 $X=587140 $Y=335740
X1136 2507 453 1 2 BUF2 $T=650380 265560 0 0 $X=650380 $Y=265180
X1137 2400 2510 1 2 BUF2 $T=651000 285720 1 0 $X=651000 $Y=280300
X1138 467 466 1 2 BUF2 $T=668360 285720 0 0 $X=668360 $Y=285340
X1139 478 2507 1 2 BUF2 $T=679520 295800 1 0 $X=679520 $Y=290380
X1140 3482 3513 1 2 BUF2 $T=1042840 315960 1 0 $X=1042840 $Y=310540
X1141 1473 1 1459 107 2 1478 ND3 $T=336040 366360 1 0 $X=336040 $Y=360940
X1142 1470 1 1436 1476 2 1478 ND3 $T=337900 356280 1 0 $X=337900 $Y=350860
X1143 1485 1 1480 1477 2 1489 ND3 $T=341620 346200 1 0 $X=341620 $Y=340780
X1144 1499 1 1476 118 2 1498 ND3 $T=346580 356280 0 0 $X=346580 $Y=355900
X1145 1499 1 122 1522 2 1505 ND3 $T=350300 356280 0 0 $X=350300 $Y=355900
X1146 1521 1 1519 1481 2 119 ND3 $T=354640 346200 0 180 $X=352160 $Y=340780
X1147 1533 1 132 123 2 129 ND3 $T=358360 366360 0 180 $X=355880 $Y=360940
X1148 145 1 1506 142 2 139 ND3 $T=364560 356280 1 180 $X=362080 $Y=355900
X1149 2019 1 2005 290 2 2013 ND3 $T=512120 356280 0 0 $X=512120 $Y=355900
X1150 2033 1 2035 296 2 2039 ND3 $T=518940 346200 0 0 $X=518940 $Y=345820
X1151 2055 1 2049 306 2 2059 ND3 $T=526380 346200 0 0 $X=526380 $Y=345820
X1152 2069 1 2065 311 2 2080 ND3 $T=529480 346200 0 0 $X=529480 $Y=345820
X1153 2051 1 2075 304 2 2081 ND3 $T=529480 356280 1 0 $X=529480 $Y=350860
X1154 2079 1 2082 310 2 2087 ND3 $T=531340 346200 1 0 $X=531340 $Y=340780
X1155 2113 1 2098 315 2 2104 ND3 $T=535680 346200 1 0 $X=535680 $Y=340780
X1156 2117 1 2121 316 2 2150 ND3 $T=540640 346200 0 0 $X=540640 $Y=345820
X1157 2138 1 2142 307 2 2159 ND3 $T=544360 356280 1 0 $X=544360 $Y=350860
X1158 330 1 2145 1955 2 329 ND3 $T=546840 366360 0 180 $X=544360 $Y=360940
X1159 2155 1 2165 331 2 2173 ND3 $T=549320 356280 1 0 $X=549320 $Y=350860
X1160 2171 1 336 337 2 2158 ND3 $T=551800 366360 0 180 $X=549320 $Y=360940
X1161 2181 1 2182 343 2 2183 ND3 $T=554280 356280 0 0 $X=554280 $Y=355900
X1162 2196 1 2176 322 2 2186 ND3 $T=554900 346200 0 0 $X=554900 $Y=345820
X1163 2189 1 2192 312 2 2197 ND3 $T=558000 336120 0 0 $X=558000 $Y=335740
X1164 2236 1 2226 355 2 2223 ND3 $T=567300 336120 0 180 $X=564820 $Y=330700
X1165 2232 1 2227 335 2 2224 ND3 $T=567300 346200 0 180 $X=564820 $Y=340780
X1166 2248 1 2252 373 2 2256 ND3 $T=572880 346200 0 0 $X=572880 $Y=345820
X1167 494 1 496 2650 2 2605 ND3 $T=701840 265560 0 0 $X=701840 $Y=265180
X1168 2631 1 489 2632 2 2618 ND3 $T=704320 305880 0 180 $X=701840 $Y=300460
X1169 499 1 496 2656 2 2646 ND3 $T=703700 265560 1 0 $X=703700 $Y=260140
X1170 2650 1 2662 491 2 2668 ND3 $T=707420 275640 1 0 $X=707420 $Y=270220
X1171 2673 1 2662 2676 2 2655 ND3 $T=709900 285720 0 180 $X=707420 $Y=280300
X1172 509 1 2684 511 2 2698 ND3 $T=714240 265560 0 0 $X=714240 $Y=265180
X1173 2653 1 2677 2703 2 2671 ND3 $T=720440 336120 0 180 $X=717960 $Y=330700
X1174 2710 1 2701 516 2 2698 ND3 $T=723540 275640 1 180 $X=721060 $Y=275260
X1175 491 1 2698 2709 2 2701 ND3 $T=721680 265560 1 0 $X=721680 $Y=260140
X1176 2691 1 2707 2714 2 2713 ND3 $T=721680 336120 1 0 $X=721680 $Y=330700
X1177 2727 1 2710 2736 2 2701 ND3 $T=733460 275640 1 180 $X=730980 $Y=275260
X1178 3072 1 3066 3046 2 3088 ND3 $T=872340 315960 0 0 $X=872340 $Y=315580
X1179 3089 1 3081 3095 2 3036 ND3 $T=880400 326040 0 180 $X=877920 $Y=320620
X1180 3255 1 3356 3342 2 3359 ND3 $T=986420 285720 1 0 $X=986420 $Y=280300
X1181 3400 1 3189 3412 2 3420 ND3 $T=1002540 305880 1 0 $X=1002540 $Y=300460
X1182 3227 1 3394 3426 2 3350 ND3 $T=1003780 315960 1 0 $X=1003780 $Y=310540
X1183 3416 1 3227 3442 2 3420 ND3 $T=1011840 305880 1 180 $X=1009360 $Y=305500
X1184 3264 1 3453 3449 2 3420 ND3 $T=1013700 315960 0 180 $X=1011220 $Y=310540
X1185 3469 1 3264 3462 2 3409 ND3 $T=1022380 305880 1 180 $X=1019900 $Y=305500
X1186 931 1 3488 3481 2 929 ND3 $T=1029200 265560 1 180 $X=1026720 $Y=265180
X1187 3508 1 941 938 2 933 ND3 $T=1032920 265560 0 180 $X=1030440 $Y=260140
X1188 3519 1 3264 3509 2 3513 ND3 $T=1036640 305880 1 180 $X=1034160 $Y=305500
X1189 995 1 986 999 2 1000 ND3 $T=1067640 265560 1 0 $X=1067640 $Y=260140
X1190 3634 1 3632 3623 2 3624 ND3 $T=1073840 285720 1 180 $X=1071360 $Y=285340
X1191 3599 1 3643 3629 2 3645 ND3 $T=1075080 315960 1 0 $X=1075080 $Y=310540
X1192 3605 1 3626 3705 2 3598 ND3 $T=1089340 295800 0 0 $X=1089340 $Y=295420
X1193 3696 1 3719 1027 2 3679 ND3 $T=1098020 285720 1 0 $X=1098020 $Y=280300
X1194 3695 1 1029 1030 2 3738 ND3 $T=1101740 265560 1 0 $X=1101740 $Y=260140
X1195 1116 1120 1122 2 1 ND2S $T=234980 275640 0 0 $X=234980 $Y=275260
X1196 90 1322 87 2 1 ND2S $T=302560 366360 0 180 $X=300700 $Y=360940
X1197 1321 1346 1325 2 1 ND2S $T=308140 336120 1 180 $X=306280 $Y=335740
X1198 1361 1351 1346 2 1 ND2S $T=311860 346200 0 180 $X=310000 $Y=340780
X1199 91 1357 1322 2 1 ND2S $T=311860 366360 0 180 $X=310000 $Y=360940
X1200 1353 1364 1349 2 1 ND2S $T=313100 346200 0 0 $X=313100 $Y=345820
X1201 1369 1303 99 2 1 ND2S $T=314960 356280 0 0 $X=314960 $Y=355900
X1202 1380 1376 99 2 1 ND2S $T=316820 336120 1 0 $X=316820 $Y=330700
X1203 1375 1345 99 2 1 ND2S $T=316820 346200 0 0 $X=316820 $Y=345820
X1204 1377 1387 1364 2 1 ND2S $T=318680 356280 1 180 $X=316820 $Y=355900
X1205 1382 1384 1308 2 1 ND2S $T=318680 326040 0 0 $X=318680 $Y=325660
X1206 1394 1397 1384 2 1 ND2S $T=321780 336120 0 180 $X=319920 $Y=330700
X1207 1391 1415 1362 2 1 ND2S $T=324260 295800 1 180 $X=322400 $Y=295420
X1208 1396 1403 1404 2 1 ND2S $T=322400 305880 0 0 $X=322400 $Y=305500
X1209 1395 1412 1355 2 1 ND2S $T=324260 315960 1 180 $X=322400 $Y=315580
X1210 1402 1411 1365 2 1 ND2S $T=325500 285720 1 180 $X=323640 $Y=285340
X1211 1413 1363 99 2 1 ND2S $T=325500 356280 1 180 $X=323640 $Y=355900
X1212 1370 1417 1407 2 1 ND2S $T=326120 275640 0 180 $X=324260 $Y=270220
X1213 1378 1443 102 2 1 ND2S $T=327360 265560 1 180 $X=325500 $Y=265180
X1214 1408 1439 1415 2 1 ND2S $T=327360 295800 1 180 $X=325500 $Y=295420
X1215 1418 1425 1403 2 1 ND2S $T=325500 305880 0 0 $X=325500 $Y=305500
X1216 1423 1428 1412 2 1 ND2S $T=327360 326040 0 180 $X=325500 $Y=320620
X1217 1424 1426 1411 2 1 ND2S $T=326740 295800 1 0 $X=326740 $Y=290380
X1218 1433 1442 1443 2 1 ND2S $T=329220 265560 0 0 $X=329220 $Y=265180
X1219 1434 1456 1417 2 1 ND2S $T=331080 275640 1 180 $X=329220 $Y=275260
X1220 1478 1469 1420 2 1 ND2S $T=338520 356280 1 180 $X=336660 $Y=355900
X1221 1478 110 1409 2 1 ND2S $T=341620 366360 0 180 $X=339760 $Y=360940
X1222 1464 1499 1507 2 1 ND2S $T=346580 336120 0 0 $X=346580 $Y=335740
X1223 1484 1505 1507 2 1 ND2S $T=350920 336120 1 180 $X=349060 $Y=335740
X1224 1514 1446 1515 2 1 ND2S $T=350920 275640 0 0 $X=350920 $Y=275260
X1225 1518 1388 1515 2 1 ND2S $T=350920 285720 1 0 $X=350920 $Y=280300
X1226 1508 1379 1515 2 1 ND2S $T=352160 305880 0 0 $X=352160 $Y=305500
X1227 1523 1393 1515 2 1 ND2S $T=354640 315960 0 180 $X=352780 $Y=310540
X1228 1517 126 1521 2 1 ND2S $T=352780 336120 1 0 $X=352780 $Y=330700
X1229 1530 1386 1515 2 1 ND2S $T=356500 305880 1 180 $X=354640 $Y=305500
X1230 1538 1416 141 2 1 ND2S $T=361460 265560 1 0 $X=361460 $Y=260140
X1231 105 1543 1552 2 1 ND2S $T=362700 295800 0 0 $X=362700 $Y=295420
X1232 1512 1645 1527 2 1 ND2S $T=388120 295800 1 0 $X=388120 $Y=290380
X1233 105 1704 1713 2 1 ND2S $T=412920 265560 0 0 $X=412920 $Y=265180
X1234 192 1541 191 2 1 ND2S $T=419740 356280 1 180 $X=417880 $Y=355900
X1235 1896 267 262 2 1 ND2S $T=482980 366360 0 180 $X=481120 $Y=360940
X1236 1933 272 1913 2 1 ND2S $T=491040 356280 1 180 $X=489180 $Y=355900
X1237 1936 1941 272 2 1 ND2S $T=492900 356280 1 180 $X=491040 $Y=355900
X1238 1949 1953 1944 2 1 ND2S $T=497860 346200 0 180 $X=496000 $Y=340780
X1239 1959 1967 1953 2 1 ND2S $T=501580 346200 0 0 $X=501580 $Y=345820
X1240 1972 1980 1962 2 1 ND2S $T=503440 346200 1 0 $X=503440 $Y=340780
X1241 1977 1995 1952 2 1 ND2S $T=510880 326040 1 180 $X=509020 $Y=325660
X1242 1996 1992 1995 2 1 ND2S $T=510880 326040 0 0 $X=510880 $Y=325660
X1243 2004 2013 2025 2 1 ND2S $T=513980 346200 1 0 $X=513980 $Y=340780
X1244 1990 2019 293 2 1 ND2S $T=514600 356280 0 0 $X=514600 $Y=355900
X1245 2017 2022 2018 2 1 ND2S $T=517700 336120 1 180 $X=515840 $Y=335740
X1246 2031 2034 2007 2 1 ND2S $T=518940 356280 1 180 $X=517080 $Y=355900
X1247 2004 2033 1989 2 1 ND2S $T=519560 346200 1 0 $X=519560 $Y=340780
X1248 2047 2039 2025 2 1 ND2S $T=521420 346200 0 0 $X=521420 $Y=345820
X1249 2048 2045 2041 2 1 ND2S $T=523900 326040 1 180 $X=522040 $Y=325660
X1250 2048 2056 2017 2 1 ND2S $T=525760 326040 1 180 $X=523900 $Y=325660
X1251 2047 2055 293 2 1 ND2S $T=526380 346200 1 180 $X=524520 $Y=345820
X1252 2066 2062 2073 2 1 ND2S $T=529480 315960 1 180 $X=527620 $Y=315580
X1253 2061 2059 2025 2 1 ND2S $T=528240 346200 1 0 $X=528240 $Y=340780
X1254 2072 2073 2076 2 1 ND2S $T=530100 315960 0 0 $X=530100 $Y=315580
X1255 2084 2081 2025 2 1 ND2S $T=533820 346200 1 180 $X=531960 $Y=345820
X1256 2061 2075 2095 2 1 ND2S $T=531960 356280 1 0 $X=531960 $Y=350860
X1257 2090 2082 2095 2 1 ND2S $T=533820 346200 1 0 $X=533820 $Y=340780
X1258 2090 2080 2025 2 1 ND2S $T=533820 346200 0 0 $X=533820 $Y=345820
X1259 2099 2096 2094 2 1 ND2S $T=536920 315960 1 180 $X=535060 $Y=315580
X1260 316 2100 314 2 1 ND2S $T=536920 356280 0 180 $X=535060 $Y=350860
X1261 2068 2094 2064 2 1 ND2S $T=537540 305880 1 180 $X=535680 $Y=305500
X1262 2084 2069 2095 2 1 ND2S $T=535680 346200 0 0 $X=535680 $Y=345820
X1263 2071 2103 2112 2 1 ND2S $T=536920 305880 1 0 $X=536920 $Y=300460
X1264 2111 2113 2095 2 1 ND2S $T=538780 346200 1 0 $X=538780 $Y=340780
X1265 2119 2128 2103 2 1 ND2S $T=542500 315960 0 180 $X=540640 $Y=310540
X1266 2111 2087 2115 2 1 ND2S $T=540640 346200 1 0 $X=540640 $Y=340780
X1267 323 319 324 2 1 ND2S $T=540640 366360 1 0 $X=540640 $Y=360940
X1268 2119 2118 2099 2 1 ND2S $T=543120 305880 0 180 $X=541260 $Y=300460
X1269 2137 2117 2095 2 1 ND2S $T=544360 336120 1 180 $X=542500 $Y=335740
X1270 307 2129 325 2 1 ND2S $T=544360 366360 0 180 $X=542500 $Y=360940
X1271 326 2136 328 2 1 ND2S $T=544360 275640 1 0 $X=544360 $Y=270220
X1272 2144 2132 2136 2 1 ND2S $T=546220 305880 1 180 $X=544360 $Y=305500
X1273 2137 2104 2115 2 1 ND2S $T=544360 346200 1 0 $X=544360 $Y=340780
X1274 2149 2138 2095 2 1 ND2S $T=546220 346200 1 180 $X=544360 $Y=345820
X1275 2149 2150 2115 2 1 ND2S $T=546840 346200 0 0 $X=546840 $Y=345820
X1276 2154 2156 2143 2 1 ND2S $T=549940 326040 0 180 $X=548080 $Y=320620
X1277 2168 2159 2115 2 1 ND2S $T=550560 346200 1 180 $X=548700 $Y=345820
X1278 2163 2167 340 2 1 ND2S $T=549940 305880 1 0 $X=549940 $Y=300460
X1279 2168 2155 2133 2 1 ND2S $T=550560 346200 0 0 $X=550560 $Y=345820
X1280 335 2105 342 2 1 ND2S $T=550560 356280 0 0 $X=550560 $Y=355900
X1281 2174 2171 325 2 1 ND2S $T=553660 366360 0 180 $X=551800 $Y=360940
X1282 2174 2152 342 2 1 ND2S $T=552420 356280 0 0 $X=552420 $Y=355900
X1283 2177 2173 2180 2 1 ND2S $T=553040 356280 1 0 $X=553040 $Y=350860
X1284 2177 2182 2133 2 1 ND2S $T=554900 356280 1 0 $X=554900 $Y=350860
X1285 2201 2186 2115 2 1 ND2S $T=558620 346200 0 180 $X=556760 $Y=340780
X1286 2190 2183 2180 2 1 ND2S $T=558000 356280 1 0 $X=558000 $Y=350860
X1287 2190 2196 2200 2 1 ND2S $T=558620 346200 0 0 $X=558620 $Y=345820
X1288 2201 2197 2200 2 1 ND2S $T=560480 346200 1 0 $X=560480 $Y=340780
X1289 2235 2174 2217 2 1 ND2S $T=562960 346200 1 0 $X=562960 $Y=340780
X1290 2213 2199 352 2 1 ND2S $T=563580 285720 0 0 $X=563580 $Y=285340
X1291 2201 2236 2169 2 1 ND2S $T=567300 326040 1 180 $X=565440 $Y=325660
X1292 2225 2223 2180 2 1 ND2S $T=565440 336120 0 0 $X=565440 $Y=335740
X1293 2218 2224 363 2 1 ND2S $T=566680 346200 0 0 $X=566680 $Y=345820
X1294 2229 2214 2233 2 1 ND2S $T=567300 305880 1 0 $X=567300 $Y=300460
X1295 2242 2192 2180 2 1 ND2S $T=570400 336120 1 180 $X=568540 $Y=335740
X1296 377 375 374 2 1 ND2S $T=577220 366360 0 180 $X=575360 $Y=360940
X1297 2212 2232 2200 2 1 ND2S $T=576600 336120 0 0 $X=576600 $Y=335740
X1298 2292 2259 386 2 1 ND2S $T=586520 295800 1 0 $X=586520 $Y=290380
X1299 2306 2294 2310 2 1 ND2S $T=590240 295800 1 0 $X=590240 $Y=290380
X1300 2308 2267 2321 2 1 ND2S $T=592720 315960 0 0 $X=592720 $Y=315580
X1301 2317 2314 2331 2 1 ND2S $T=593340 326040 0 0 $X=593340 $Y=325660
X1302 2331 2303 2330 2 1 ND2S $T=595200 326040 0 0 $X=595200 $Y=325660
X1303 2323 2302 2336 2 1 ND2S $T=595820 315960 0 0 $X=595820 $Y=315580
X1304 2350 2280 2373 2 1 ND2S $T=608220 336120 0 0 $X=608220 $Y=335740
X1305 2379 2322 2383 2 1 ND2S $T=610080 346200 1 0 $X=610080 $Y=340780
X1306 2385 2304 2378 2 1 ND2S $T=611940 356280 0 0 $X=611940 $Y=355900
X1307 2392 2290 2374 2 1 ND2S $T=615040 326040 0 0 $X=615040 $Y=325660
X1308 2417 2359 2407 2 1 ND2S $T=620620 356280 0 0 $X=620620 $Y=355900
X1309 2587 2590 2603 2 1 ND2S $T=686340 275640 1 0 $X=686340 $Y=270220
X1310 2592 2609 2587 2 1 ND2S $T=693780 275640 1 180 $X=691920 $Y=275260
X1311 487 485 491 2 1 ND2S $T=693160 265560 1 0 $X=693160 $Y=260140
X1312 2623 2614 2629 2 1 ND2S $T=698740 285720 1 0 $X=698740 $Y=280300
X1313 2617 2638 2664 2 1 ND2S $T=703700 295800 1 0 $X=703700 $Y=290380
X1314 2640 2641 2631 2 1 ND2S $T=706180 285720 0 0 $X=706180 $Y=285340
X1315 2666 2665 2627 2 1 ND2S $T=708040 305880 1 180 $X=706180 $Y=305500
X1316 2627 2652 2670 2 1 ND2S $T=708040 305880 1 0 $X=708040 $Y=300460
X1317 2666 2662 2631 2 1 ND2S $T=708660 295800 0 0 $X=708660 $Y=295420
X1318 2671 2648 2677 2 1 ND2S $T=709280 326040 0 0 $X=709280 $Y=325660
X1319 2680 2668 506 2 1 ND2S $T=714240 275640 0 180 $X=712380 $Y=270220
X1320 512 2695 2682 2 1 ND2S $T=717960 336120 0 0 $X=717960 $Y=335740
X1321 2715 512 518 2 1 ND2S $T=721680 346200 1 0 $X=721680 $Y=340780
X1322 518 2730 2740 2 1 ND2S $T=734080 356280 1 0 $X=734080 $Y=350860
X1323 2739 2747 2727 2 1 ND2S $T=739660 275640 1 180 $X=737800 $Y=275260
X1324 518 2753 2749 2 1 ND2S $T=740900 326040 0 180 $X=739040 $Y=320620
X1325 2698 2762 2739 2 1 ND2S $T=745240 285720 0 180 $X=743380 $Y=280300
X1326 2765 2789 2728 2 1 ND2S $T=753300 326040 0 180 $X=751440 $Y=320620
X1327 2765 2807 2798 2 1 ND2S $T=757020 326040 0 180 $X=755160 $Y=320620
X1328 2765 2839 2776 2 1 ND2S $T=770040 315960 1 180 $X=768180 $Y=315580
X1329 2765 2849 2834 2 1 ND2S $T=771900 326040 0 180 $X=770040 $Y=320620
X1330 2765 2862 2840 2 1 ND2S $T=776860 336120 0 180 $X=775000 $Y=330700
X1331 2765 2857 2818 2 1 ND2S $T=776860 336120 1 180 $X=775000 $Y=335740
X1332 2715 2878 2881 2 1 ND2S $T=781820 346200 1 0 $X=781820 $Y=340780
X1333 2877 2881 2857 2 1 ND2S $T=784300 346200 1 0 $X=784300 $Y=340780
X1334 596 2893 2903 2 1 ND2S $T=789260 275640 1 0 $X=789260 $Y=270220
X1335 2911 592 593 2 1 ND2S $T=794220 265560 1 0 $X=794220 $Y=260140
X1336 2911 2918 606 2 1 ND2S $T=803520 265560 1 0 $X=803520 $Y=260140
X1337 2911 2944 609 2 1 ND2S $T=809100 265560 0 180 $X=807240 $Y=260140
X1338 606 618 621 2 1 ND2S $T=811580 265560 1 0 $X=811580 $Y=260140
X1339 2957 2950 606 2 1 ND2S $T=812820 265560 0 0 $X=812820 $Y=265180
X1340 2957 2921 593 2 1 ND2S $T=813440 265560 1 0 $X=813440 $Y=260140
X1341 619 2968 2963 2 1 ND2S $T=817780 285720 1 0 $X=817780 $Y=280300
X1342 2911 2969 2903 2 1 ND2S $T=820880 265560 1 0 $X=820880 $Y=260140
X1343 2957 2967 609 2 1 ND2S $T=823980 265560 1 0 $X=823980 $Y=260140
X1344 624 2986 2989 2 1 ND2S $T=828320 285720 0 180 $X=826460 $Y=280300
X1345 648 2987 2984 2 1 ND2S $T=828320 305880 0 180 $X=826460 $Y=300460
X1346 2957 2992 2903 2 1 ND2S $T=830180 265560 0 180 $X=828320 $Y=260140
X1347 2976 2988 2999 2 1 ND2S $T=830180 346200 1 0 $X=830180 $Y=340780
X1348 660 2995 606 2 1 ND2S $T=833900 285720 1 0 $X=833900 $Y=280300
X1349 2911 3000 2963 2 1 ND2S $T=835760 265560 0 0 $X=835760 $Y=265180
X1350 2957 3015 2963 2 1 ND2S $T=841960 265560 1 180 $X=840100 $Y=265180
X1351 2911 3017 2989 2 1 ND2S $T=843820 265560 0 0 $X=843820 $Y=265180
X1352 705 3008 593 2 1 ND2S $T=858700 285720 0 0 $X=858700 $Y=285340
X1353 3082 3069 2989 2 1 ND2S $T=872340 265560 0 0 $X=872340 $Y=265180
X1354 717 3074 720 2 1 ND2S $T=876680 265560 0 0 $X=876680 $Y=265180
X1355 3066 3105 3081 2 1 ND2S $T=877920 315960 0 0 $X=877920 $Y=315580
X1356 840 3309 3266 2 1 ND2S $T=969060 285720 0 180 $X=967200 $Y=280300
X1357 840 3307 3235 2 1 ND2S $T=969060 295800 0 180 $X=967200 $Y=290380
X1358 840 3316 3255 2 1 ND2S $T=972780 275640 1 180 $X=970920 $Y=275260
X1359 846 3301 3235 2 1 ND2S $T=972160 285720 1 0 $X=972160 $Y=280300
X1360 846 3306 3189 2 1 ND2S $T=972780 295800 0 0 $X=972780 $Y=295420
X1361 846 3314 3266 2 1 ND2S $T=974020 275640 0 0 $X=974020 $Y=275260
X1362 3350 3335 774 2 1 ND2S $T=982700 265560 1 0 $X=982700 $Y=260140
X1363 846 863 3255 2 1 ND2S $T=985180 275640 1 180 $X=983320 $Y=275260
X1364 3357 871 3361 2 1 ND2S $T=987040 366360 1 0 $X=987040 $Y=360940
X1365 3350 3392 3227 2 1 ND2S $T=997580 315960 0 180 $X=995720 $Y=310540
X1366 3395 887 3398 2 1 ND2S $T=996340 366360 1 0 $X=996340 $Y=360940
X1367 803 3323 3411 2 1 ND2S $T=1000680 265560 0 0 $X=1000680 $Y=265180
X1368 888 3427 892 2 1 ND2S $T=1006260 275640 0 180 $X=1004400 $Y=270220
X1369 3420 3425 803 2 1 ND2S $T=1007500 265560 1 180 $X=1005640 $Y=265180
X1370 3450 906 3434 2 1 ND2S $T=1009980 265560 1 180 $X=1008120 $Y=265180
X1371 3425 3434 3445 2 1 ND2S $T=1008120 275640 1 0 $X=1008120 $Y=270220
X1372 3229 3445 3350 2 1 ND2S $T=1011220 275640 1 0 $X=1011220 $Y=270220
X1373 3449 3444 3454 2 1 ND2S $T=1011220 326040 1 0 $X=1011220 $Y=320620
X1374 3229 911 3359 2 1 ND2S $T=1013080 275640 1 0 $X=1013080 $Y=270220
X1375 3429 3454 3457 2 1 ND2S $T=1013080 315960 0 0 $X=1013080 $Y=315580
X1376 3350 3489 3264 2 1 ND2S $T=1023620 305880 0 0 $X=1023620 $Y=305500
X1377 3227 3480 3482 2 1 ND2S $T=1023620 315960 1 0 $X=1023620 $Y=310540
X1378 3411 3500 3189 2 1 ND2S $T=1027960 315960 0 180 $X=1026100 $Y=310540
X1379 3359 3494 3281 2 1 ND2S $T=1031060 305880 0 180 $X=1029200 $Y=300460
X1380 3281 3497 3411 2 1 ND2S $T=1031060 315960 0 180 $X=1029200 $Y=310540
X1381 3501 3495 3493 2 1 ND2S $T=1031060 326040 1 180 $X=1029200 $Y=325660
X1382 3515 3496 3518 2 1 ND2S $T=1034780 275640 1 0 $X=1034780 $Y=270220
X1383 3507 3519 3492 2 1 ND2S $T=1037880 305880 0 0 $X=1037880 $Y=305500
X1384 3506 941 972 2 1 ND2S $T=1045320 265560 0 0 $X=1045320 $Y=265180
X1385 983 3523 991 2 1 ND2S $T=1054620 265560 1 0 $X=1054620 $Y=260140
X1386 3484 3550 3565 2 1 ND2S $T=1055860 315960 0 0 $X=1055860 $Y=315580
X1387 3569 3565 3571 2 1 ND2S $T=1057720 326040 1 180 $X=1055860 $Y=325660
X1388 989 3532 3566 2 1 ND2S $T=1058340 275640 0 180 $X=1056480 $Y=270220
X1389 3559 3590 3576 2 1 ND2S $T=1061440 305880 0 180 $X=1059580 $Y=300460
X1390 3577 3569 3568 2 1 ND2S $T=1059580 326040 0 0 $X=1059580 $Y=325660
X1391 3484 3588 3576 2 1 ND2S $T=1062060 295800 1 180 $X=1060200 $Y=295420
X1392 3590 3578 3596 2 1 ND2S $T=1062680 315960 1 0 $X=1062680 $Y=310540
X1393 3589 3592 3584 2 1 ND2S $T=1063300 326040 0 0 $X=1063300 $Y=325660
X1394 3608 3583 3614 2 1 ND2S $T=1068260 285720 0 0 $X=1068260 $Y=285340
X1395 3609 3604 3614 2 1 ND2S $T=1068260 295800 1 0 $X=1068260 $Y=290380
X1396 3618 3585 3625 2 1 ND2S $T=1070120 275640 0 0 $X=1070120 $Y=275260
X1397 3635 3602 3617 2 1 ND2S $T=1073840 326040 0 0 $X=1073840 $Y=325660
X1398 3596 3651 3652 2 1 ND2S $T=1076940 315960 0 0 $X=1076940 $Y=315580
X1399 3650 3663 3629 2 1 ND2S $T=1081280 305880 0 180 $X=1079420 $Y=300460
X1400 3607 3639 3680 2 1 ND2S $T=1084380 295800 0 0 $X=1084380 $Y=295420
X1401 3659 3622 3667 2 1 ND2S $T=1084380 326040 0 0 $X=1084380 $Y=325660
X1402 3636 3677 3626 2 1 ND2S $T=1087480 305880 1 0 $X=1087480 $Y=300460
X1403 3689 3696 3707 2 1 ND2S $T=1093680 275640 0 0 $X=1093680 $Y=275260
X1404 3710 3723 3697 2 1 ND2S $T=1098640 265560 1 180 $X=1096780 $Y=265180
X1405 3718 3700 3751 2 1 ND2S $T=1099880 326040 0 0 $X=1099880 $Y=325660
X1406 3718 3720 3698 2 1 ND2S $T=1104220 326040 1 180 $X=1102360 $Y=325660
X1407 3724 3739 3726 2 1 ND2S $T=1106080 275640 1 180 $X=1104220 $Y=275260
X1408 3734 3735 3747 2 1 ND2S $T=1104220 315960 0 0 $X=1104220 $Y=315580
X1409 3753 3734 3756 2 1 ND2S $T=1106700 315960 0 0 $X=1106700 $Y=315580
X1410 3752 3714 3754 2 1 ND2S $T=1107320 275640 0 0 $X=1107320 $Y=275260
X1411 3755 3751 3741 2 1 ND2S $T=1107320 326040 1 0 $X=1107320 $Y=320620
X1412 3770 3775 3762 2 1 ND2S $T=1112280 326040 0 180 $X=1110420 $Y=320620
X1413 3765 3770 3741 2 1 ND2S $T=1111040 336120 1 0 $X=1111040 $Y=330700
X1414 3773 3763 3776 2 1 ND2S $T=1112280 295800 0 0 $X=1112280 $Y=295420
X1415 1043 1041 1040 2 1 ND2S $T=1114760 265560 0 180 $X=1112900 $Y=260140
X1416 3761 3769 3754 2 1 ND2S $T=1114760 285720 1 0 $X=1114760 $Y=280300
X1417 3798 1043 3797 2 1 ND2S $T=1119720 265560 1 0 $X=1119720 $Y=260140
X1418 3761 3799 3797 2 1 ND2S $T=1125300 265560 0 0 $X=1125300 $Y=265180
X1419 1086 6 1 5 1077 1074 2 MOAI1S $T=224440 285720 1 180 $X=220720 $Y=285340
X1420 1093 6 1 10 9 1079 2 MOAI1S $T=225680 265560 1 180 $X=221960 $Y=265180
X1421 1099 16 1 5 1085 1081 2 MOAI1S $T=226920 346200 1 180 $X=223200 $Y=345820
X1422 1084 1091 1 5 1096 1080 2 MOAI1S $T=223820 305880 1 0 $X=223820 $Y=300460
X1423 1098 16 1 5 1092 1076 2 MOAI1S $T=227540 315960 1 180 $X=223820 $Y=315580
X1424 23 6 1 10 24 1078 2 MOAI1S $T=233740 265560 1 0 $X=233740 $Y=260140
X1425 133 1512 1 1534 1537 1529 2 MOAI1S $T=357120 295800 1 0 $X=357120 $Y=290380
X1426 133 1539 1 138 1543 1500 2 MOAI1S $T=359600 305880 1 0 $X=359600 $Y=300460
X1427 174 1697 1 186 1704 189 2 MOAI1S $T=408580 265560 1 0 $X=408580 $Y=260140
X1428 2592 2584 1 2592 2590 2572 2 MOAI1S $T=686960 275640 1 180 $X=683240 $Y=275260
X1429 2600 2615 1 2609 2614 2616 2 MOAI1S $T=695020 285720 1 0 $X=695020 $Y=280300
X1430 495 497 1 495 497 2660 2 MOAI1S $T=701840 356280 0 0 $X=701840 $Y=355900
X1431 482 500 1 2637 2654 2658 2 MOAI1S $T=703700 275640 1 0 $X=703700 $Y=270220
X1432 2653 2661 1 2653 2648 2644 2 MOAI1S $T=708660 326040 1 180 $X=704940 $Y=325660
X1433 2667 2663 1 2667 2663 2657 2 MOAI1S $T=711140 356280 1 180 $X=707420 $Y=355900
X1434 2670 2665 1 2666 2638 2679 2 MOAI1S $T=709280 305880 0 0 $X=709280 $Y=305500
X1435 2684 500 1 2684 2654 2699 2 MOAI1S $T=714860 275640 1 0 $X=714860 $Y=270220
X1436 519 2717 1 519 2709 523 2 MOAI1S $T=724780 265560 1 0 $X=724780 $Y=260140
X1437 2639 2706 1 2714 2705 2697 2 MOAI1S $T=724780 315960 0 0 $X=724780 $Y=315580
X1438 2701 2712 1 2687 2727 2723 2 MOAI1S $T=727260 275640 0 0 $X=727260 $Y=275260
X1439 2707 2724 1 2707 2703 2718 2 MOAI1S $T=732220 326040 1 180 $X=728500 $Y=325660
X1440 524 2726 1 524 2726 2732 2 MOAI1S $T=729120 265560 1 0 $X=729120 $Y=260140
X1441 2689 2730 1 2689 2730 2737 2 MOAI1S $T=731600 326040 1 0 $X=731600 $Y=320620
X1442 527 2732 1 527 2732 2764 2 MOAI1S $T=733460 265560 1 0 $X=733460 $Y=260140
X1443 2742 2731 1 2742 2741 2725 2 MOAI1S $T=738420 315960 0 180 $X=734700 $Y=310540
X1444 2734 2753 1 2734 2753 2752 2 MOAI1S $T=744000 315960 1 180 $X=740280 $Y=315580
X1445 2754 2761 1 2754 2761 2759 2 MOAI1S $T=744620 315960 0 180 $X=740900 $Y=310540
X1446 2774 2772 1 2774 2772 2769 2 MOAI1S $T=748960 315960 0 180 $X=745240 $Y=310540
X1447 2782 2789 1 2782 2789 2799 2 MOAI1S $T=749580 315960 1 0 $X=749580 $Y=310540
X1448 2771 2764 1 2771 2764 2813 2 MOAI1S $T=753300 275640 1 0 $X=753300 $Y=270220
X1449 2802 2807 1 2802 2807 2816 2 MOAI1S $T=755780 315960 0 0 $X=755780 $Y=315580
X1450 2817 2820 1 2817 2820 2814 2 MOAI1S $T=763840 315960 0 180 $X=760120 $Y=310540
X1451 2831 2839 1 2831 2839 2835 2 MOAI1S $T=770660 315960 0 180 $X=766940 $Y=310540
X1452 2847 2849 1 2847 2849 2855 2 MOAI1S $T=771280 315960 0 0 $X=771280 $Y=315580
X1453 2828 2864 1 2828 2864 2871 2 MOAI1S $T=778100 315960 0 0 $X=778100 $Y=315580
X1454 2859 2862 1 2859 2862 2875 2 MOAI1S $T=778100 336120 1 0 $X=778100 $Y=330700
X1455 2882 2874 1 2762 577 2854 2 MOAI1S $T=783060 305880 1 180 $X=779340 $Y=305500
X1456 2858 2872 1 2858 2883 2899 2 MOAI1S $T=782440 326040 1 0 $X=782440 $Y=320620
X1457 2880 2884 1 2880 2889 2900 2 MOAI1S $T=783060 326040 0 0 $X=783060 $Y=325660
X1458 2762 2897 1 2762 581 2888 2 MOAI1S $T=789260 305880 1 180 $X=785540 $Y=305500
X1459 2904 2898 1 2904 2898 2919 2 MOAI1S $T=796080 346200 1 0 $X=796080 $Y=340780
X1460 2882 2941 1 2882 604 2932 2 MOAI1S $T=805380 315960 1 180 $X=801660 $Y=315580
X1461 2882 2956 1 2882 614 2938 2 MOAI1S $T=813440 315960 1 180 $X=809720 $Y=315580
X1462 2960 2913 1 2960 2913 2949 2 MOAI1S $T=819640 346200 0 180 $X=815920 $Y=340780
X1463 2971 2975 1 2971 632 2966 2 MOAI1S $T=823360 315960 1 180 $X=819640 $Y=315580
X1464 634 2968 1 634 2968 2965 2 MOAI1S $T=824600 285720 0 180 $X=820880 $Y=280300
X1465 2971 2978 1 2971 643 2983 2 MOAI1S $T=822740 315960 1 0 $X=822740 $Y=310540
X1466 2991 2987 1 2991 2987 2998 2 MOAI1S $T=828320 305880 1 0 $X=828320 $Y=300460
X1467 2986 2995 1 2986 2995 2974 2 MOAI1S $T=833900 285720 0 180 $X=830180 $Y=280300
X1468 3003 2988 1 3003 2988 2996 2 MOAI1S $T=833900 346200 1 0 $X=833900 $Y=340780
X1469 2971 3010 1 3014 674 3022 2 MOAI1S $T=840720 315960 1 0 $X=840720 $Y=310540
X1470 2738 3047 1 3036 3054 3045 2 MOAI1S $T=858700 326040 1 0 $X=858700 $Y=320620
X1471 3014 3050 1 3014 703 3053 2 MOAI1S $T=864280 305880 0 180 $X=860560 $Y=300460
X1472 3014 3070 1 3014 711 3064 2 MOAI1S $T=869240 295800 1 180 $X=865520 $Y=295420
X1473 3066 3072 1 3066 3072 3020 2 MOAI1S $T=871100 326040 0 180 $X=867380 $Y=320620
X1474 3083 3095 1 3083 3095 3110 2 MOAI1S $T=876060 326040 0 0 $X=876060 $Y=325660
X1475 3099 3106 1 3099 722 3098 2 MOAI1S $T=882260 285720 0 180 $X=878540 $Y=280300
X1476 3099 3111 1 3099 729 3113 2 MOAI1S $T=881640 295800 0 0 $X=881640 $Y=295420
X1477 3089 3105 1 3089 3105 3120 2 MOAI1S $T=881640 315960 0 0 $X=881640 $Y=315580
X1478 3099 3148 1 3099 742 3153 2 MOAI1S $T=899620 285720 1 0 $X=899620 $Y=280300
X1479 3158 3167 1 3158 577 3142 2 MOAI1S $T=910780 305880 0 180 $X=907060 $Y=300460
X1480 752 3175 1 2736 674 3161 2 MOAI1S $T=912640 275640 1 180 $X=908920 $Y=275260
X1481 3174 3155 1 3174 632 3162 2 MOAI1S $T=913260 326040 1 180 $X=909540 $Y=325660
X1482 3158 3181 1 3158 614 3168 2 MOAI1S $T=914500 295800 1 180 $X=910780 $Y=295420
X1483 3180 3177 1 3180 581 3141 2 MOAI1S $T=915740 315960 0 180 $X=912020 $Y=310540
X1484 752 755 1 752 703 3182 2 MOAI1S $T=917600 275640 0 180 $X=913880 $Y=270220
X1485 3174 3144 1 3174 604 3179 2 MOAI1S $T=923180 326040 1 180 $X=919460 $Y=325660
X1486 3203 3212 1 3203 770 769 2 MOAI1S $T=928760 356280 1 180 $X=925040 $Y=355900
X1487 3174 3222 1 3174 643 3211 2 MOAI1S $T=931240 336120 0 180 $X=927520 $Y=330700
X1488 777 779 1 777 742 773 2 MOAI1S $T=931860 265560 1 180 $X=928140 $Y=265180
X1489 2747 3223 1 2747 703 3192 2 MOAI1S $T=931860 275640 1 180 $X=928140 $Y=275260
X1490 3218 3224 1 3218 577 3207 2 MOAI1S $T=931860 305880 0 180 $X=928140 $Y=300460
X1491 758 3219 1 758 770 3214 2 MOAI1S $T=932480 356280 1 180 $X=928760 $Y=355900
X1492 758 3183 1 758 781 3231 2 MOAI1S $T=930000 346200 1 0 $X=930000 $Y=340780
X1493 3218 3230 1 3218 581 3216 2 MOAI1S $T=934960 305880 1 180 $X=931240 $Y=305500
X1494 2747 3232 1 2747 722 3226 2 MOAI1S $T=935580 275640 1 180 $X=931860 $Y=275260
X1495 3218 3220 1 3218 604 3225 2 MOAI1S $T=938680 315960 0 180 $X=934960 $Y=310540
X1496 3203 790 1 3203 786 3228 2 MOAI1S $T=938680 366360 0 180 $X=934960 $Y=360940
X1497 3203 3246 1 3203 781 3252 2 MOAI1S $T=941780 346200 0 0 $X=941780 $Y=345820
X1498 3253 3256 1 3253 674 3245 2 MOAI1S $T=948600 275640 1 180 $X=944880 $Y=275260
X1499 3254 3257 1 3254 643 3244 2 MOAI1S $T=948600 315960 1 180 $X=944880 $Y=315580
X1500 3253 3258 1 3253 614 3247 2 MOAI1S $T=949220 295800 1 180 $X=945500 $Y=295420
X1501 3253 3265 1 791 742 3241 2 MOAI1S $T=952940 265560 1 180 $X=949220 $Y=265180
X1502 3254 3267 1 3254 632 3260 2 MOAI1S $T=952940 315960 1 180 $X=949220 $Y=315580
X1503 806 3275 1 806 781 3280 2 MOAI1S $T=954800 346200 0 0 $X=954800 $Y=345820
X1504 726 3271 1 806 3286 3287 2 MOAI1S $T=959140 346200 0 0 $X=959140 $Y=345820
X1505 3145 3298 1 3291 781 3290 2 MOAI1S $T=966580 346200 1 180 $X=962860 $Y=345820
X1506 3291 3313 1 3291 839 3292 2 MOAI1S $T=970920 356280 1 180 $X=967200 $Y=355900
X1507 3291 3315 1 3291 3286 3320 2 MOAI1S $T=970300 346200 0 0 $X=970300 $Y=345820
X1508 3329 3328 1 3329 3328 3288 2 MOAI1S $T=980840 275640 1 180 $X=977120 $Y=275260
X1509 859 3353 1 859 857 3334 2 MOAI1S $T=983940 366360 0 180 $X=980220 $Y=360940
X1510 3356 3355 1 3356 3355 3328 2 MOAI1S $T=989520 275640 1 180 $X=985800 $Y=275260
X1511 3369 3377 1 3369 857 3333 2 MOAI1S $T=993860 356280 0 180 $X=990140 $Y=350860
X1512 859 3384 1 859 885 3388 2 MOAI1S $T=992620 366360 1 0 $X=992620 $Y=360940
X1513 3394 3392 1 3394 3392 3375 2 MOAI1S $T=998820 305880 1 180 $X=995100 $Y=305500
X1514 3402 3400 1 3402 3400 3336 2 MOAI1S $T=1001300 305880 0 180 $X=997580 $Y=300460
X1515 3419 3416 1 3419 3416 3408 2 MOAI1S $T=1006880 305880 1 180 $X=1003160 $Y=305500
X1516 3413 3369 1 3369 885 3415 2 MOAI1S $T=1003160 346200 0 0 $X=1003160 $Y=345820
X1517 898 3424 1 898 885 896 2 MOAI1S $T=1006880 366360 0 180 $X=1003160 $Y=360940
X1518 903 3440 1 903 885 3433 2 MOAI1S $T=1011220 356280 0 180 $X=1007500 $Y=350860
X1519 3436 3435 1 888 3448 3450 2 MOAI1S $T=1008740 275640 0 0 $X=1008740 $Y=275260
X1520 903 3455 1 903 857 3463 2 MOAI1S $T=1013080 356280 1 0 $X=1013080 $Y=350860
X1521 898 3459 1 898 857 916 2 MOAI1S $T=1014940 366360 1 0 $X=1014940 $Y=360940
X1522 3453 3461 1 3453 3461 3460 2 MOAI1S $T=1016180 315960 1 0 $X=1016180 $Y=310540
X1523 3460 3462 1 3460 3462 3466 2 MOAI1S $T=1016180 315960 0 0 $X=1016180 $Y=315580
X1524 3469 3464 1 3469 3464 3431 2 MOAI1S $T=1021760 305880 0 180 $X=1018040 $Y=300460
X1525 3369 3467 1 3369 917 3472 2 MOAI1S $T=1018040 356280 1 0 $X=1018040 $Y=350860
X1526 898 3476 1 898 917 3470 2 MOAI1S $T=1023000 366360 0 180 $X=1019280 $Y=360940
X1527 3405 3479 1 3405 3479 3483 2 MOAI1S $T=1021760 336120 1 0 $X=1021760 $Y=330700
X1528 932 3496 1 3499 942 3505 2 MOAI1S $T=1029200 275640 1 0 $X=1029200 $Y=270220
X1529 3511 3509 1 3511 3509 3498 2 MOAI1S $T=1036640 336120 0 180 $X=1032920 $Y=330700
X1530 3510 3514 1 3510 917 3520 2 MOAI1S $T=1033540 356280 1 0 $X=1033540 $Y=350860
X1531 3528 949 1 3518 3521 3512 2 MOAI1S $T=1040980 275640 0 180 $X=1037260 $Y=270220
X1532 3522 3483 1 3522 3483 3511 2 MOAI1S $T=1040980 336120 0 180 $X=1037260 $Y=330700
X1533 3525 3497 1 3525 3497 3522 2 MOAI1S $T=1042220 315960 1 180 $X=1038500 $Y=315580
X1534 964 3539 1 3541 3539 3542 2 MOAI1S $T=1045940 275640 0 0 $X=1045940 $Y=275260
X1535 3549 3552 1 3549 917 3546 2 MOAI1S $T=1050280 356280 1 0 $X=1050280 $Y=350860
X1536 3484 3582 1 3578 3573 3556 2 MOAI1S $T=1062680 315960 0 180 $X=1058960 $Y=310540
X1537 3543 3583 1 3543 3583 3593 2 MOAI1S $T=1060820 285720 0 0 $X=1060820 $Y=285340
X1538 993 3585 1 993 3585 3579 2 MOAI1S $T=1065160 265560 1 180 $X=1061440 $Y=265180
X1539 3570 3604 1 3570 3604 3600 2 MOAI1S $T=1070120 285720 0 180 $X=1066400 $Y=280300
X1540 3592 3595 1 3592 3595 3615 2 MOAI1S $T=1066400 336120 1 0 $X=1066400 $Y=330700
X1541 3626 3603 1 3613 3602 3610 2 MOAI1S $T=1071980 315960 0 180 $X=1068260 $Y=310540
X1542 1003 3601 1 1003 1002 3508 2 MOAI1S $T=1074460 265560 0 180 $X=1070740 $Y=260140
X1543 3631 1003 1 3631 1003 3644 2 MOAI1S $T=1072600 275640 0 0 $X=1072600 $Y=275260
X1544 3635 3617 1 3635 3617 3641 2 MOAI1S $T=1073220 336120 1 0 $X=1073220 $Y=330700
X1545 3655 3633 1 3655 3632 3625 2 MOAI1S $T=1081900 285720 0 180 $X=1078180 $Y=280300
X1546 3596 3657 1 3651 3666 3658 2 MOAI1S $T=1078800 315960 0 0 $X=1078800 $Y=315580
X1547 3656 1009 1 3656 1009 3670 2 MOAI1S $T=1079420 265560 1 0 $X=1079420 $Y=260140
X1548 3655 3663 1 3655 3647 3609 2 MOAI1S $T=1083140 295800 0 180 $X=1079420 $Y=290380
X1549 3647 3655 1 3663 3638 3679 2 MOAI1S $T=1081900 285720 0 0 $X=1081900 $Y=285340
X1550 3638 3647 1 3638 3633 3662 2 MOAI1S $T=1086240 285720 0 180 $X=1082520 $Y=280300
X1551 3636 3628 1 3677 3598 3684 2 MOAI1S $T=1083760 305880 1 0 $X=1083760 $Y=300460
X1552 3690 3666 1 3605 3681 3669 2 MOAI1S $T=1090580 315960 0 180 $X=1086860 $Y=310540
X1553 3686 3691 1 3696 3649 3701 2 MOAI1S $T=1089340 275640 0 0 $X=1089340 $Y=275260
X1554 3706 3697 1 3695 1022 3673 2 MOAI1S $T=1093680 265560 0 180 $X=1089960 $Y=260140
X1555 3729 3726 1 3719 3649 3745 2 MOAI1S $T=1101740 285720 1 0 $X=1101740 $Y=280300
X1556 3705 3746 1 3705 3746 3736 2 MOAI1S $T=1107940 295800 0 180 $X=1104220 $Y=290380
X1557 3759 1034 1 1029 1022 3740 2 MOAI1S $T=1109180 265560 0 180 $X=1105460 $Y=260140
X1558 3761 3758 1 3769 3752 3777 2 MOAI1S $T=1109800 285720 1 0 $X=1109800 $Y=280300
X1559 3774 3750 1 3774 3750 3781 2 MOAI1S $T=1111660 315960 1 0 $X=1111660 $Y=310540
X1560 3765 3741 1 3765 3741 3784 2 MOAI1S $T=1119100 326040 1 180 $X=1115380 $Y=325660
X1561 3763 3787 1 3763 3787 3796 2 MOAI1S $T=1123440 295800 1 180 $X=1119720 $Y=295420
X1562 3761 3766 1 3799 3798 3792 2 MOAI1S $T=1125300 265560 1 180 $X=1121580 $Y=265180
X1563 1349 2 1352 1353 1 NR2 $T=314960 346200 0 180 $X=313100 $Y=340780
X1564 1308 2 1401 1382 1 NR2 $T=320540 326040 0 180 $X=318680 $Y=320620
X1565 1365 2 1421 1402 1 NR2 $T=321780 285720 0 0 $X=321780 $Y=285340
X1566 1404 2 1405 1396 1 NR2 $T=324260 305880 0 180 $X=322400 $Y=300460
X1567 102 2 1429 1378 1 NR2 $T=326120 265560 1 0 $X=326120 $Y=260140
X1568 1409 2 1459 1420 1 NR2 $T=336660 356280 1 180 $X=334800 $Y=355900
X1569 1462 2 1473 1436 1 NR2 $T=337900 356280 0 180 $X=336040 $Y=350860
X1570 1477 2 1478 1481 1 NR2 $T=339760 346200 0 0 $X=339760 $Y=345820
X1571 1480 2 1488 1481 1 NR2 $T=341620 346200 0 0 $X=341620 $Y=345820
X1572 1486 2 114 1482 1 NR2 $T=341620 356280 0 0 $X=341620 $Y=355900
X1573 1448 2 1489 1484 1 NR2 $T=342240 336120 0 0 $X=342240 $Y=335740
X1574 1488 2 1498 1496 1 NR2 $T=348440 346200 0 180 $X=346580 $Y=340780
X1575 1448 2 1507 1481 1 NR2 $T=348440 346200 1 0 $X=348440 $Y=340780
X1576 121 2 1502 1504 1 NR2 $T=350920 326040 0 180 $X=349060 $Y=320620
X1577 121 2 1513 1520 1 NR2 $T=351540 326040 1 0 $X=351540 $Y=320620
X1578 131 2 119 137 1 NR2 $T=355880 346200 1 0 $X=355880 $Y=340780
X1579 1533 2 1525 1526 1 NR2 $T=357740 356280 1 0 $X=357740 $Y=350860
X1580 140 2 1533 144 1 NR2 $T=362700 356280 1 0 $X=362700 $Y=350860
X1581 1570 2 143 142 1 NR2 $T=364560 366360 0 180 $X=362700 $Y=360940
X1582 154 2 1589 1624 1 NR2 $T=386260 295800 1 0 $X=386260 $Y=290380
X1583 1626 2 1609 1607 1 NR2 $T=388120 326040 0 180 $X=386260 $Y=320620
X1584 153 2 1631 1632 1 NR2 $T=387500 275640 1 0 $X=387500 $Y=270220
X1585 155 2 1616 154 1 NR2 $T=389360 285720 0 180 $X=387500 $Y=280300
X1586 1626 2 1629 1628 1 NR2 $T=388120 326040 0 0 $X=388120 $Y=325660
X1587 157 2 1597 1632 1 NR2 $T=389360 275640 1 0 $X=389360 $Y=270220
X1588 161 2 1605 154 1 NR2 $T=391220 285720 0 180 $X=389360 $Y=280300
X1589 1643 2 1627 1628 1 NR2 $T=391220 336120 1 180 $X=389360 $Y=335740
X1590 162 2 1630 1637 1 NR2 $T=391220 356280 0 180 $X=389360 $Y=350860
X1591 160 2 156 164 1 NR2 $T=389980 356280 0 0 $X=389980 $Y=355900
X1592 1607 2 1608 1649 1 NR2 $T=390600 305880 1 0 $X=390600 $Y=300460
X1593 162 2 1638 165 1 NR2 $T=390600 326040 0 0 $X=390600 $Y=325660
X1594 1645 2 168 138 1 NR2 $T=391220 285720 0 0 $X=391220 $Y=285340
X1595 1637 2 1594 1619 1 NR2 $T=391220 295800 1 0 $X=391220 $Y=290380
X1596 1653 2 1598 1619 1 NR2 $T=393080 326040 0 180 $X=391220 $Y=320620
X1597 1650 2 1646 1628 1 NR2 $T=393080 346200 1 180 $X=391220 $Y=345820
X1598 163 2 1636 1628 1 NR2 $T=391220 356280 1 0 $X=391220 $Y=350860
X1599 154 2 1651 1619 1 NR2 $T=391840 275640 0 0 $X=391840 $Y=275260
X1600 155 2 1633 1649 1 NR2 $T=391840 285720 1 0 $X=391840 $Y=280300
X1601 1650 2 1610 165 1 NR2 $T=391840 346200 1 0 $X=391840 $Y=340780
X1602 153 2 167 1624 1 NR2 $T=392460 265560 1 0 $X=392460 $Y=260140
X1603 1637 2 1642 1652 1 NR2 $T=394320 305880 0 180 $X=392460 $Y=300460
X1604 163 2 1614 1655 1 NR2 $T=392460 326040 0 0 $X=392460 $Y=325660
X1605 169 2 1621 166 1 NR2 $T=394940 356280 1 180 $X=393080 $Y=355900
X1606 1643 2 1639 166 1 NR2 $T=393700 356280 1 0 $X=393700 $Y=350860
X1607 1626 2 1640 1657 1 NR2 $T=394320 295800 1 0 $X=394320 $Y=290380
X1608 1643 2 1661 1660 1 NR2 $T=394320 305880 0 0 $X=394320 $Y=305500
X1609 1659 2 1654 163 1 NR2 $T=396180 326040 1 180 $X=394320 $Y=325660
X1610 157 2 1648 1624 1 NR2 $T=394940 265560 1 0 $X=394940 $Y=260140
X1611 170 2 1613 1649 1 NR2 $T=396800 275640 1 180 $X=394940 $Y=275260
X1612 157 2 1656 1649 1 NR2 $T=396800 285720 0 180 $X=394940 $Y=280300
X1613 170 2 1634 1643 1 NR2 $T=396800 295800 1 180 $X=394940 $Y=295420
X1614 1660 2 1625 1649 1 NR2 $T=396800 305880 0 180 $X=394940 $Y=300460
X1615 1643 2 1664 1668 1 NR2 $T=394940 326040 1 0 $X=394940 $Y=320620
X1616 163 2 1635 1668 1 NR2 $T=394940 336120 1 0 $X=394940 $Y=330700
X1617 163 2 1663 165 1 NR2 $T=394940 336120 0 0 $X=394940 $Y=335740
X1618 1650 2 1665 1655 1 NR2 $T=398660 326040 1 180 $X=396800 $Y=325660
X1619 1653 2 1673 164 1 NR2 $T=396800 336120 0 0 $X=396800 $Y=335740
X1620 1653 2 1641 1657 1 NR2 $T=399280 295800 0 180 $X=397420 $Y=290380
X1621 1643 2 1670 1655 1 NR2 $T=397420 305880 0 0 $X=397420 $Y=305500
X1622 1607 2 1674 1637 1 NR2 $T=398660 305880 1 0 $X=398660 $Y=300460
X1623 1653 2 1667 1668 1 NR2 $T=398660 326040 1 0 $X=398660 $Y=320620
X1624 1659 2 1669 1650 1 NR2 $T=400520 326040 1 180 $X=398660 $Y=325660
X1625 1650 2 1676 1668 1 NR2 $T=398660 336120 1 0 $X=398660 $Y=330700
X1626 1619 2 1675 1649 1 NR2 $T=401760 295800 0 180 $X=399900 $Y=290380
X1627 176 2 1666 1677 1 NR2 $T=399900 346200 0 0 $X=399900 $Y=345820
X1628 1653 2 1678 1607 1 NR2 $T=401140 326040 0 0 $X=401140 $Y=325660
X1629 181 2 1679 1624 1 NR2 $T=403620 265560 0 180 $X=401760 $Y=260140
X1630 161 2 1683 1632 1 NR2 $T=403620 285720 0 180 $X=401760 $Y=280300
X1631 1619 2 1698 1624 1 NR2 $T=402380 285720 0 0 $X=402380 $Y=285340
X1632 1626 2 1681 1668 1 NR2 $T=404240 326040 0 180 $X=402380 $Y=320620
X1633 1637 2 1690 180 1 NR2 $T=402380 346200 0 0 $X=402380 $Y=345820
X1634 179 2 1680 180 1 NR2 $T=402380 366360 1 0 $X=402380 $Y=360940
X1635 181 2 1684 1632 1 NR2 $T=403620 265560 1 0 $X=403620 $Y=260140
X1636 1626 2 1699 165 1 NR2 $T=405480 305880 1 180 $X=403620 $Y=305500
X1637 1652 2 1685 180 1 NR2 $T=405480 315960 0 180 $X=403620 $Y=310540
X1638 161 2 1702 1624 1 NR2 $T=404240 265560 0 0 $X=404240 $Y=265180
X1639 1691 2 1692 165 1 NR2 $T=406100 356280 0 180 $X=404240 $Y=350860
X1640 170 2 1687 1653 1 NR2 $T=406720 295800 0 180 $X=404860 $Y=290380
X1641 179 2 1695 1652 1 NR2 $T=407340 326040 0 180 $X=405480 $Y=320620
X1642 1691 2 1689 1655 1 NR2 $T=407340 336120 0 180 $X=405480 $Y=330700
X1643 179 2 1696 175 1 NR2 $T=407340 366360 0 180 $X=405480 $Y=360940
X1644 183 2 1686 1691 1 NR2 $T=409820 326040 1 180 $X=407960 $Y=325660
X1645 170 2 1705 179 1 NR2 $T=409200 285720 0 0 $X=409200 $Y=285340
X1646 188 2 1703 1677 1 NR2 $T=411680 356280 0 180 $X=409820 $Y=350860
X1647 183 2 1707 188 1 NR2 $T=412300 356280 1 0 $X=412300 $Y=350860
X1648 188 2 1706 184 1 NR2 $T=414780 356280 1 180 $X=412920 $Y=355900
X1649 192 2 1712 1731 1 NR2 $T=418500 346200 1 0 $X=418500 $Y=340780
X1650 198 2 1506 195 1 NR2 $T=422840 356280 1 180 $X=420980 $Y=355900
X1651 199 2 1570 201 1 NR2 $T=423460 366360 1 0 $X=423460 $Y=360940
X1652 145 2 1752 1731 1 NR2 $T=429660 346200 0 0 $X=429660 $Y=345820
X1653 217 2 1756 1731 1 NR2 $T=433380 346200 1 180 $X=431520 $Y=345820
X1654 1772 2 1753 1731 1 NR2 $T=434000 356280 0 180 $X=432140 $Y=350860
X1655 209 2 1765 1731 1 NR2 $T=435240 346200 1 180 $X=433380 $Y=345820
X1656 220 2 1773 219 1 NR2 $T=436480 366360 0 180 $X=434620 $Y=360940
X1657 262 2 263 1896 1 NR2 $T=479260 366360 1 0 $X=479260 $Y=360940
X1658 1913 2 271 1933 1 NR2 $T=488560 366360 1 0 $X=488560 $Y=360940
X1659 1944 2 1956 1949 1 NR2 $T=496620 336120 0 0 $X=496620 $Y=335740
X1660 1929 2 1969 1965 1 NR2 $T=499720 336120 1 0 $X=499720 $Y=330700
X1661 1969 2 1973 1974 1 NR2 $T=502820 336120 1 0 $X=502820 $Y=330700
X1662 1952 2 1974 1977 1 NR2 $T=506540 326040 0 0 $X=506540 $Y=325660
X1663 318 2 2109 2114 1 NR2 $T=538160 356280 1 0 $X=538160 $Y=350860
X1664 318 2 2139 2091 1 NR2 $T=544360 356280 1 180 $X=542500 $Y=355900
X1665 2140 2 2131 327 1 NR2 $T=545600 305880 0 180 $X=543740 $Y=300460
X1666 362 2 2228 360 1 NR2 $T=569160 275640 0 180 $X=567300 $Y=270220
X1667 371 2 368 209 1 NR2 $T=572260 366360 0 180 $X=570400 $Y=360940
X1668 371 2 2258 1772 1 NR2 $T=575980 356280 1 180 $X=574120 $Y=355900
X1669 379 2 2268 2264 1 NR2 $T=580940 295800 1 180 $X=579080 $Y=295420
X1670 371 2 2293 384 1 NR2 $T=587760 346200 1 0 $X=587760 $Y=340780
X1671 392 2 393 394 1 NR2 $T=589000 366360 1 0 $X=589000 $Y=360940
X1672 2311 2 2317 2329 1 NR2 $T=595820 326040 1 0 $X=595820 $Y=320620
X1673 2341 2 2311 2348 1 NR2 $T=598920 305880 1 0 $X=598920 $Y=300460
X1674 2368 2 2360 2364 1 NR2 $T=607600 315960 1 180 $X=605740 $Y=315580
X1675 2365 2 2335 2370 1 NR2 $T=606360 346200 0 0 $X=606360 $Y=345820
X1676 2376 2 2355 2390 1 NR2 $T=611940 346200 1 0 $X=611940 $Y=340780
X1677 2398 2 2384 2365 1 NR2 $T=616280 356280 1 180 $X=614420 $Y=355900
X1678 2402 2 2390 2394 1 NR2 $T=616280 336120 0 0 $X=616280 $Y=335740
X1679 2415 2 2376 2410 1 NR2 $T=620620 346200 0 180 $X=618760 $Y=340780
X1680 2441 2 2365 2434 1 NR2 $T=627440 356280 0 0 $X=627440 $Y=355900
X1681 426 2 2398 2447 1 NR2 $T=633020 356280 1 180 $X=631160 $Y=355900
X1682 2295 2 2459 422 1 NR2 $T=635500 356280 1 180 $X=633640 $Y=355900
X1683 2618 2 2627 489 1 NR2 $T=699360 305880 1 180 $X=697500 $Y=305500
X1684 2622 2 2629 2625 1 NR2 $T=698740 275640 0 0 $X=698740 $Y=275260
X1685 2627 2 2626 2631 1 NR2 $T=699980 305880 1 0 $X=699980 $Y=300460
X1686 493 2 2634 489 1 NR2 $T=700600 305880 0 0 $X=700600 $Y=305500
X1687 2625 2 2605 2633 1 NR2 $T=703700 275640 1 180 $X=701840 $Y=275260
X1688 2634 2 2666 2638 1 NR2 $T=702460 305880 0 0 $X=702460 $Y=305500
X1689 2632 2 2651 2640 1 NR2 $T=705560 305880 1 0 $X=705560 $Y=300460
X1690 498 2 2667 2660 1 NR2 $T=706180 366360 1 0 $X=706180 $Y=360940
X1691 502 2 2646 2662 1 NR2 $T=707420 265560 0 0 $X=707420 $Y=265180
X1692 509 2 507 2656 1 NR2 $T=714860 265560 0 180 $X=713000 $Y=260140
X1693 2659 2 2681 2671 1 NR2 $T=713000 326040 0 0 $X=713000 $Y=325660
X1694 2690 2 2687 500 1 NR2 $T=717960 275640 1 180 $X=716100 $Y=275260
X1695 2701 2 2690 2654 1 NR2 $T=720440 275640 1 180 $X=718580 $Y=275260
X1696 512 2 2671 2691 1 NR2 $T=718580 346200 1 0 $X=718580 $Y=340780
X1697 2698 2 2712 2654 1 NR2 $T=721680 275640 0 180 $X=719820 $Y=270220
X1698 2677 2 2713 2653 1 NR2 $T=723540 336120 0 0 $X=723540 $Y=335740
X1699 2704 2 2739 521 1 NR2 $T=734700 275640 0 180 $X=732840 $Y=270220
X1700 2705 2 2742 2737 1 NR2 $T=736560 315960 1 180 $X=734700 $Y=315580
X1701 2705 2 2754 2752 1 NR2 $T=737800 315960 0 0 $X=737800 $Y=315580
X1702 2773 2 2774 2799 1 NR2 $T=755780 315960 0 180 $X=753920 $Y=310540
X1703 2773 2 2817 2816 1 NR2 $T=757640 315960 1 0 $X=757640 $Y=310540
X1704 2773 2 2828 2835 1 NR2 $T=764460 315960 1 0 $X=764460 $Y=310540
X1705 2838 2 2858 2855 1 NR2 $T=777480 315960 1 180 $X=775620 $Y=315580
X1706 2838 2 2880 2875 1 NR2 $T=780580 326040 0 0 $X=780580 $Y=325660
X1707 2877 2 2902 2857 1 NR2 $T=788020 346200 0 180 $X=786160 $Y=340780
X1708 2918 2 2908 2921 1 NR2 $T=797320 265560 1 0 $X=797320 $Y=260140
X1709 2944 2 2930 2950 1 NR2 $T=809100 265560 1 0 $X=809100 $Y=260140
X1710 2969 2 2959 2967 1 NR2 $T=821500 265560 0 0 $X=821500 $Y=265180
X1711 651 2 2991 649 1 NR2 $T=830180 285720 0 180 $X=828320 $Y=280300
X1712 3000 2 653 2992 1 NR2 $T=832040 265560 0 180 $X=830180 $Y=260140
X1713 3017 2 3016 3015 1 NR2 $T=843820 265560 1 180 $X=841960 $Y=265180
X1714 3056 2 3047 3036 1 NR2 $T=862420 326040 1 0 $X=862420 $Y=320620
X1715 3056 2 3025 3063 1 NR2 $T=864280 326040 0 0 $X=864280 $Y=325660
X1716 3056 2 3066 3063 1 NR2 $T=864900 326040 1 0 $X=864900 $Y=320620
X1717 3074 2 3055 3069 1 NR2 $T=869860 265560 0 0 $X=869860 $Y=265180
X1718 3083 2 3088 3089 1 NR2 $T=874820 315960 0 0 $X=874820 $Y=315580
X1719 3309 2 3299 3301 1 NR2 $T=969060 275640 0 0 $X=969060 $Y=275260
X1720 3307 2 3305 3306 1 NR2 $T=970920 295800 0 0 $X=970920 $Y=295420
X1721 3316 2 3289 3314 1 NR2 $T=973400 265560 1 0 $X=973400 $Y=260140
X1722 3335 2 3294 3323 1 NR2 $T=978980 265560 1 0 $X=978980 $Y=260140
X1723 3354 2 3337 3346 1 NR2 $T=983320 285720 1 180 $X=981460 $Y=285340
X1724 3354 2 3341 3351 1 NR2 $T=984560 285720 0 180 $X=982700 $Y=280300
X1725 3342 2 3331 3336 1 NR2 $T=982700 295800 0 0 $X=982700 $Y=295420
X1726 3354 2 3303 3322 1 NR2 $T=983320 285720 0 0 $X=983320 $Y=285340
X1727 873 2 3330 3368 1 NR2 $T=988280 285720 0 0 $X=988280 $Y=285340
X1728 877 2 3355 3351 1 NR2 $T=992000 285720 0 180 $X=990140 $Y=280300
X1729 877 2 3358 3366 1 NR2 $T=993860 275640 0 180 $X=992000 $Y=270220
X1730 882 2 3356 3366 1 NR2 $T=993860 285720 0 180 $X=992000 $Y=280300
X1731 3368 2 3381 3351 1 NR2 $T=992000 285720 0 0 $X=992000 $Y=285340
X1732 3370 2 3376 3375 1 NR2 $T=992000 315960 1 0 $X=992000 $Y=310540
X1733 3382 2 3371 3376 1 NR2 $T=993860 326040 0 180 $X=992000 $Y=320620
X1734 873 2 3380 3354 1 NR2 $T=993860 265560 0 0 $X=993860 $Y=265180
X1735 873 2 3378 882 1 NR2 $T=993860 275640 1 0 $X=993860 $Y=270220
X1736 882 2 3393 3351 1 NR2 $T=995720 285720 0 180 $X=993860 $Y=280300
X1737 3389 2 3386 3366 1 NR2 $T=995720 285720 1 180 $X=993860 $Y=285340
X1738 888 2 3373 3389 1 NR2 $T=997580 275640 0 180 $X=995720 $Y=270220
X1739 3396 2 3391 3346 1 NR2 $T=997580 285720 1 180 $X=995720 $Y=285340
X1740 3396 2 3374 3322 1 NR2 $T=996960 285720 1 0 $X=996960 $Y=280300
X1741 888 2 3399 877 1 NR2 $T=997580 265560 0 0 $X=997580 $Y=265180
X1742 892 2 3401 3389 1 NR2 $T=1000680 275640 0 180 $X=998820 $Y=270220
X1743 3368 2 3404 3322 1 NR2 $T=1000680 285720 1 180 $X=998820 $Y=285340
X1744 3410 2 3385 3322 1 NR2 $T=1001300 285720 0 180 $X=999440 $Y=280300
X1745 3412 2 3403 3408 1 NR2 $T=1002540 305880 1 180 $X=1000680 $Y=305500
X1746 888 2 899 3354 1 NR2 $T=1004400 265560 1 0 $X=1004400 $Y=260140
X1747 3410 2 3422 3346 1 NR2 $T=1006260 285720 1 180 $X=1004400 $Y=285340
X1748 3396 2 3428 3438 1 NR2 $T=1007500 285720 0 0 $X=1007500 $Y=285340
X1749 3430 2 3402 3438 1 NR2 $T=1007500 305880 1 0 $X=1007500 $Y=300460
X1750 3430 2 3419 3439 1 NR2 $T=1007500 305880 0 0 $X=1007500 $Y=305500
X1751 3410 2 3443 3438 1 NR2 $T=1009360 285720 0 0 $X=1009360 $Y=285340
X1752 3368 2 3446 3346 1 NR2 $T=1011840 285720 0 180 $X=1009980 $Y=280300
X1753 3436 2 3390 3438 1 NR2 $T=1009980 295800 1 0 $X=1009980 $Y=290380
X1754 3448 2 3400 3439 1 NR2 $T=1011840 305880 0 180 $X=1009980 $Y=300460
X1755 3442 2 3429 3431 1 NR2 $T=1009980 315960 0 0 $X=1009980 $Y=315580
X1756 3439 2 3451 3368 1 NR2 $T=1013080 285720 1 180 $X=1011220 $Y=285340
X1757 3396 2 3473 3439 1 NR2 $T=1014940 285720 1 180 $X=1013080 $Y=285340
X1758 3436 2 3453 3456 1 NR2 $T=1013080 295800 1 0 $X=1013080 $Y=290380
X1759 3448 2 3416 3456 1 NR2 $T=1013080 305880 1 0 $X=1013080 $Y=300460
X1760 3430 2 3461 3458 1 NR2 $T=1014940 305880 1 0 $X=1014940 $Y=300460
X1761 3396 2 3468 3458 1 NR2 $T=1015560 295800 1 0 $X=1015560 $Y=290380
X1762 3448 2 3464 3458 1 NR2 $T=1016800 295800 0 0 $X=1016800 $Y=295420
X1763 3430 2 3469 3456 1 NR2 $T=1018660 295800 0 0 $X=1018660 $Y=295420
X1764 3460 2 3478 3462 1 NR2 $T=1022380 315960 0 180 $X=1020520 $Y=310540
X1765 3456 2 3477 3410 1 NR2 $T=1021760 295800 0 0 $X=1021760 $Y=295420
X1766 3466 2 3471 3426 1 NR2 $T=1023000 326040 1 0 $X=1023000 $Y=320620
X1767 3489 2 3492 3494 1 NR2 $T=1032300 305880 0 0 $X=1032300 $Y=305500
X1768 3506 2 3499 3512 1 NR2 $T=1032920 275640 1 0 $X=1032920 $Y=270220
X1769 3480 2 3507 3500 1 NR2 $T=1036020 315960 1 0 $X=1036020 $Y=310540
X1770 963 2 965 3528 1 NR2 $T=1043460 265560 1 0 $X=1043460 $Y=260140
X1771 3528 2 939 975 1 NR2 $T=1045320 265560 1 0 $X=1045320 $Y=260140
X1772 3547 2 3517 3542 1 NR2 $T=1050280 285720 1 180 $X=1048420 $Y=285340
X1773 3559 2 3533 3558 1 NR2 $T=1057100 315960 0 180 $X=1055240 $Y=310540
X1774 983 2 990 991 1 NR2 $T=1059580 265560 0 180 $X=1057720 $Y=260140
X1775 3569 2 3559 3571 1 NR2 $T=1057720 326040 1 0 $X=1057720 $Y=320620
X1776 3547 2 3564 3579 1 NR2 $T=1058960 275640 1 0 $X=1058960 $Y=270220
X1777 3567 2 3582 3590 1 NR2 $T=1059580 315960 0 0 $X=1059580 $Y=315580
X1778 3547 2 3587 3593 1 NR2 $T=1065160 295800 0 180 $X=1063300 $Y=290380
X1779 3547 2 3594 3600 1 NR2 $T=1064540 285720 1 0 $X=1064540 $Y=280300
X1780 3590 2 3598 3573 1 NR2 $T=1067020 305880 1 180 $X=1065160 $Y=305500
X1781 3605 2 3603 3590 1 NR2 $T=1068260 315960 0 180 $X=1066400 $Y=310540
X1782 3582 2 3607 3610 1 NR2 $T=1067640 305880 0 0 $X=1067640 $Y=305500
X1783 3615 2 3536 3627 1 NR2 $T=1070120 336120 1 0 $X=1070120 $Y=330700
X1784 3634 2 3630 3639 1 NR2 $T=1073840 295800 1 0 $X=1073840 $Y=290380
X1785 3642 2 3618 3646 1 NR2 $T=1075700 285720 1 0 $X=1075700 $Y=280300
X1786 3634 2 3642 3645 1 NR2 $T=1075700 305880 1 0 $X=1075700 $Y=300460
X1787 3649 2 3653 3644 1 NR2 $T=1078800 275640 1 180 $X=1076940 $Y=275260
X1788 3629 2 3647 3619 1 NR2 $T=1079420 295800 0 180 $X=1077560 $Y=290380
X1789 3654 2 3664 3627 1 NR2 $T=1078800 336120 1 0 $X=1078800 $Y=330700
X1790 3642 2 3656 3662 1 NR2 $T=1079420 275640 0 0 $X=1079420 $Y=275260
X1791 3649 2 1017 3670 1 NR2 $T=1085000 265560 0 180 $X=1083140 $Y=260140
X1792 3626 2 3628 3681 1 NR2 $T=1084380 315960 1 0 $X=1084380 $Y=310540
X1793 3652 2 3657 3678 1 NR2 $T=1084380 315960 0 0 $X=1084380 $Y=315580
X1794 3689 2 3686 3547 1 NR2 $T=1089340 275640 1 180 $X=1087480 $Y=275260
X1795 3710 2 3706 1024 1 NR2 $T=1094920 265560 1 0 $X=1094920 $Y=260140
X1796 3714 2 3710 3707 1 NR2 $T=1096780 275640 0 180 $X=1094920 $Y=270220
X1797 3724 2 3729 3649 1 NR2 $T=1103600 275640 0 180 $X=1101740 $Y=270220
X1798 3736 2 3712 3732 1 NR2 $T=1103600 295800 1 180 $X=1101740 $Y=295420
X1799 3734 2 3666 3747 1 NR2 $T=1102360 305880 0 0 $X=1102360 $Y=305500
X1800 3698 2 3760 3627 1 NR2 $T=1107320 336120 1 0 $X=1107320 $Y=330700
X1801 3705 2 3773 3746 1 NR2 $T=1111040 295800 1 180 $X=1109180 $Y=295420
X1802 1036 2 3759 1022 1 NR2 $T=1109800 265560 1 0 $X=1109800 $Y=260140
X1803 3770 2 3753 3762 1 NR2 $T=1112900 315960 0 0 $X=1112900 $Y=315580
X1804 3785 2 3786 3627 1 NR2 $T=1116000 336120 0 180 $X=1114140 $Y=330700
X1805 3763 2 3752 3787 1 NR2 $T=1114760 295800 0 0 $X=1114760 $Y=295420
X1806 3788 2 3793 3732 1 NR2 $T=1116000 305880 0 0 $X=1116000 $Y=305500
X1807 3795 2 3789 3732 1 NR2 $T=1119100 295800 1 180 $X=1117240 $Y=295420
X1808 3797 2 3766 3739 1 NR2 $T=1121580 265560 1 180 $X=1119720 $Y=265180
X1809 2848 480 1 2 INV12CK $T=771900 366360 0 180 $X=761980 $Y=360940
X1810 2848 557 1 2 INV12CK $T=784920 356280 0 0 $X=784920 $Y=355900
X1811 3149 669 1 2 INV12CK $T=900240 366360 0 180 $X=890320 $Y=360940
X1812 3149 659 1 2 INV12CK $T=904580 326040 0 180 $X=894660 $Y=320620
X1813 865 905 1 2 INV12CK $T=1006260 356280 0 0 $X=1006260 $Y=355900
X1814 1195 67 2 1 1243 OR2 $T=269700 336120 0 0 $X=269700 $Y=335740
X1815 1186 1218 2 1 1262 OR2 $T=279000 295800 0 0 $X=279000 $Y=295420
X1816 1321 1325 2 1 1361 OR2 $T=305660 346200 1 0 $X=305660 $Y=340780
X1817 1391 1362 2 1 1408 OR2 $T=321780 295800 1 0 $X=321780 $Y=290380
X1818 1395 1355 2 1 1423 OR2 $T=321780 326040 1 0 $X=321780 $Y=320620
X1819 1370 1407 2 1 1434 OR2 $T=326120 275640 1 0 $X=326120 $Y=270220
X1820 1501 1488 2 1 124 OR2 $T=348440 356280 1 0 $X=348440 $Y=350860
X1821 1504 125 2 1 128 OR2 $T=352160 315960 0 0 $X=352160 $Y=315580
X1822 1731 192 2 1 1719 OR2 $T=420360 356280 0 180 $X=417880 $Y=350860
X1823 1721 1719 2 1 1730 OR2 $T=419740 275640 1 0 $X=419740 $Y=270220
X1824 2028 2020 2 1 2017 OR2 $T=517080 326040 1 180 $X=514600 $Y=325660
X1825 2038 2011 2 1 2048 OR2 $T=522660 315960 1 0 $X=522660 $Y=310540
X1826 2072 2076 2 1 2066 OR2 $T=531960 315960 0 180 $X=529480 $Y=310540
X1827 2068 2064 2 1 2099 OR2 $T=535060 315960 1 0 $X=535060 $Y=310540
X1828 2071 2112 2 1 2119 OR2 $T=538780 305880 0 0 $X=538780 $Y=305500
X1829 326 328 2 1 2144 OR2 $T=543740 275640 0 0 $X=543740 $Y=275260
X1830 192 371 2 1 374 OR2 $T=572260 366360 1 0 $X=572260 $Y=360940
X1831 2382 2249 2 1 2396 OR2 $T=613180 315960 0 0 $X=613180 $Y=315580
X1832 2481 2482 2 1 2494 OR2 $T=641700 315960 0 0 $X=641700 $Y=315580
X1833 518 2705 2 1 2706 OR2 $T=724160 315960 1 180 $X=721680 $Y=315580
X1834 2878 2902 2 1 2904 OR2 $T=789260 346200 1 0 $X=789260 $Y=340780
X1835 3068 3056 2 1 3078 OR2 $T=867380 326040 0 0 $X=867380 $Y=325660
X1836 3194 2680 2 1 3202 OR2 $T=920700 295800 1 0 $X=920700 $Y=290380
X1837 3194 3484 2 1 3502 OR2 $T=1025480 295800 0 0 $X=1025480 $Y=295420
X1838 3650 3629 2 1 3633 OR2 $T=1078800 305880 0 0 $X=1078800 $Y=305500
X1839 3726 3723 2 1 3719 OR2 $T=1100500 275640 1 180 $X=1098020 $Y=275260
X1840 2636 2640 2641 2630 2 1 2655 OA22 $T=702460 285720 1 0 $X=702460 $Y=280300
X1841 1101 1089 1 2 1105 AN2 $T=227540 336120 1 0 $X=227540 $Y=330700
X1842 1217 1126 1 2 1209 AN2 $T=265980 295800 0 180 $X=263500 $Y=290380
X1843 75 79 1 2 1265 AN2 $T=280860 366360 1 0 $X=280860 $Y=360940
X1844 81 79 1 2 1274 AN2 $T=284580 366360 1 0 $X=284580 $Y=360940
X1845 1285 79 1 2 1291 AN2 $T=290780 346200 0 0 $X=290780 $Y=345820
X1846 1269 79 1 2 1290 AN2 $T=291400 336120 1 0 $X=291400 $Y=330700
X1847 1289 1316 1 2 1320 AN2 $T=300700 315960 1 0 $X=300700 $Y=310540
X1848 1312 1316 1 2 1323 AN2 $T=301940 285720 0 0 $X=301940 $Y=285340
X1849 1331 1316 1 2 1340 AN2 $T=305660 305880 1 0 $X=305660 $Y=300460
X1850 1311 79 1 2 1343 AN2 $T=305660 315960 0 0 $X=305660 $Y=315580
X1851 1298 95 1 2 1359 AN2 $T=307520 265560 0 0 $X=307520 $Y=265180
X1852 1297 1316 1 2 96 AN2 $T=309380 265560 1 0 $X=309380 $Y=260140
X1853 1327 1316 1 2 1354 AN2 $T=309380 275640 1 0 $X=309380 $Y=270220
X1854 2220 366 1 2 2246 AN2 $T=568540 336120 1 0 $X=568540 $Y=330700
X1855 501 498 1 2 2659 AN2 $T=704320 336120 0 0 $X=704320 $Y=335740
X1856 3370 3375 1 2 3382 AN2 $T=991380 305880 0 0 $X=991380 $Y=305500
X1857 3409 3427 1 2 3435 AN2 $T=1005640 275640 0 0 $X=1005640 $Y=275260
X1858 3634 3647 1 2 3646 AN2 $T=1077560 285720 0 0 $X=1077560 $Y=285340
X1859 3666 3652 1 2 3659 AN2 $T=1087480 326040 1 0 $X=1087480 $Y=320620
X1860 3598 3626 1 2 3699 AN2 $T=1089340 305880 1 0 $X=1089340 $Y=300460
X1861 1522 2 1525 124 134 1 NR3 $T=354020 356280 0 0 $X=354020 $Y=355900
X1862 2620 2 2664 2631 2680 1 NR3 $T=714240 295800 1 180 $X=711140 $Y=295420
X1863 3628 2 3657 3669 3645 1 NR3 $T=1080040 315960 1 0 $X=1080040 $Y=310540
X1864 3758 2 3766 3772 3738 1 NR3 $T=1109800 275640 0 0 $X=1109800 $Y=275260
X1865 31 1149 1 1152 2 OR2B1S $T=243040 346200 1 0 $X=243040 $Y=340780
X1866 31 1140 1 1161 2 OR2B1S $T=243660 326040 0 0 $X=243660 $Y=325660
X1867 1154 1114 1 1168 2 OR2B1S $T=248620 285720 1 0 $X=248620 $Y=280300
X1868 1154 49 1 1185 2 OR2B1S $T=257920 265560 1 180 $X=254820 $Y=265180
X1869 1159 1196 1 1239 2 OR2B1S $T=268460 305880 0 0 $X=268460 $Y=305500
X1870 1901 1902 1 1909 2 OR2B1S $T=480500 336120 1 0 $X=480500 $Y=330700
X1871 1987 2161 1 2146 2 OR2B1S $T=554280 295800 1 180 $X=551180 $Y=295420
X1872 2239 2205 1 2234 2 OR2B1S $T=569780 315960 1 180 $X=566680 $Y=315580
X1873 2239 2016 1 2261 2 OR2B1S $T=574120 326040 1 0 $X=574120 $Y=320620
X1874 2239 2257 1 2273 2 OR2B1S $T=578460 285720 1 0 $X=578460 $Y=280300
X1875 2445 2454 1 2485 2 OR2B1S $T=634260 326040 0 0 $X=634260 $Y=325660
X1876 2445 2462 1 2478 2 OR2B1S $T=636740 346200 1 0 $X=636740 $Y=340780
X1877 2239 442 1 2500 2 OR2B1S $T=644800 315960 0 0 $X=644800 $Y=315580
X1878 2638 2626 1 2625 2 OR2B1S $T=702460 285720 1 180 $X=699360 $Y=285340
X1879 506 2680 1 2673 2 OR2B1S $T=712380 275640 0 0 $X=712380 $Y=275260
X1880 2712 2687 1 2717 2 OR2B1S $T=724160 275640 0 0 $X=724160 $Y=275260
X1881 2733 2673 1 2722 2 OR2B1S $T=734080 295800 1 180 $X=730980 $Y=295420
X1882 3576 3559 1 3597 2 OR2B1S $T=1062060 305880 0 0 $X=1062060 $Y=305500
X1883 3697 3710 1 3695 2 OR2B1S $T=1096780 265560 1 0 $X=1096780 $Y=260140
X1884 637 2848 1 2 INV6CK $T=822740 356280 0 0 $X=822740 $Y=355900
X1885 637 3149 1 2 INV6CK $T=903960 356280 0 0 $X=903960 $Y=355900
X1886 637 865 1 2 INV6CK $T=982080 356280 0 0 $X=982080 $Y=355900
X1887 1965 1962 1929 1 2 ND2 $T=501580 336120 1 180 $X=499720 $Y=335740
X1888 2028 2018 2020 1 2 ND2 $T=517080 326040 0 0 $X=517080 $Y=325660
X1889 2038 2041 2011 1 2 ND2 $T=523280 315960 0 0 $X=523280 $Y=315580
X1890 327 2143 2140 1 2 ND2 $T=545600 305880 1 0 $X=545600 $Y=300460
X1891 334 2158 324 1 2 ND2 $T=549320 366360 0 180 $X=547460 $Y=360940
X1892 2144 2170 2154 1 2 ND2 $T=551180 315960 0 180 $X=549320 $Y=310540
X1893 360 2233 362 1 2 ND2 $T=566680 275640 0 0 $X=566680 $Y=275260
X1894 2212 2256 363 1 2 ND2 $T=575360 346200 0 0 $X=575360 $Y=345820
X1895 2225 2252 2200 1 2 ND2 $T=577220 346200 0 0 $X=577220 $Y=345820
X1896 2320 2310 399 1 2 ND2 $T=593960 285720 1 0 $X=593960 $Y=280300
X1897 2333 2336 2342 1 2 ND2 $T=597680 315960 1 0 $X=597680 $Y=310540
X1898 2339 2345 2335 1 2 ND2 $T=599540 356280 0 180 $X=597680 $Y=350860
X1899 2339 2334 2350 1 2 ND2 $T=599540 336120 0 0 $X=599540 $Y=335740
X1900 2339 2344 2355 1 2 ND2 $T=599540 346200 1 0 $X=599540 $Y=340780
X1901 2348 2321 2341 1 2 ND2 $T=601400 305880 1 0 $X=601400 $Y=300460
X1902 2364 2330 2368 1 2 ND2 $T=606360 315960 1 0 $X=606360 $Y=310540
X1903 2394 2373 2402 1 2 ND2 $T=614420 336120 0 0 $X=614420 $Y=335740
X1904 2395 2374 2401 1 2 ND2 $T=615040 326040 1 0 $X=615040 $Y=320620
X1905 2410 2383 2415 1 2 ND2 $T=618760 346200 0 0 $X=618760 $Y=345820
X1906 2434 2378 2441 1 2 ND2 $T=625580 356280 0 0 $X=625580 $Y=355900
X1907 2447 2407 426 1 2 ND2 $T=629300 366360 1 0 $X=629300 $Y=360940
X1908 1469 1476 1506 123 2 1 127 OA112 $T=347820 366360 1 0 $X=347820 $Y=360940
X1909 313 308 2091 2092 2 1 317 OA112 $T=533200 366360 1 0 $X=533200 $Y=360940
X1910 3596 3592 3589 3584 2 1 3580 OA112 $T=1065160 336120 0 180 $X=1060200 $Y=330700
X1911 3596 3622 3659 3667 2 1 3674 OA112 $T=1078180 326040 0 0 $X=1078180 $Y=325660
X1912 3636 3705 3699 3708 2 1 3716 OA112 $T=1092440 295800 0 0 $X=1092440 $Y=295420
X1913 3636 3720 3718 3698 2 1 3711 OA112 $T=1099880 326040 1 180 $X=1094920 $Y=325660
X1914 3636 3763 3773 3776 2 1 3767 OA112 $T=1109180 305880 1 0 $X=1109180 $Y=300460
X1915 2625 2622 1 2641 500 2617 2 OAI112HS $T=703700 275640 0 0 $X=703700 $Y=275260
X1916 3633 3630 1 3623 3539 3618 2 OAI112HS $T=1074460 285720 0 180 $X=1070120 $Y=280300
X1917 333 2 2170 1 2184 NR2P $T=554900 315960 1 0 $X=554900 $Y=310540
X1918 2228 2 357 1 2240 NR2P $T=569780 285720 1 180 $X=566060 $Y=285340
X1919 2301 2 379 1 2260 NR2P $T=587760 285720 0 0 $X=587760 $Y=285340
X1920 399 2 2320 1 2301 NR2P $T=595820 285720 1 0 $X=595820 $Y=280300
X1921 2342 2 2333 1 2329 NR2P $T=599540 315960 1 0 $X=599540 $Y=310540
X1922 2363 2 2360 1 2347 NR2P $T=603260 326040 0 0 $X=603260 $Y=325660
X1923 2401 2 2395 1 2363 NR2P $T=616900 326040 1 0 $X=616900 $Y=320620
X1924 111 110 1469 2 1490 1 113 AN4B1S $T=341620 366360 1 0 $X=341620 $Y=360940
X1925 2100 2052 2105 2 2109 1 320 AN4B1S $T=536300 356280 0 0 $X=536300 $Y=355900
X1926 2129 2078 2152 2 2139 1 2145 AN4B1S $T=546220 356280 0 0 $X=546220 $Y=355900
X1927 3597 3620 3607 2 3628 1 3616 AN4B1S $T=1069500 305880 0 0 $X=1069500 $Y=305500
X1928 3597 3614 3645 2 3582 1 3650 AN4B1S $T=1074460 305880 0 0 $X=1074460 $Y=305500
X1929 1118 2 28 1104 32 1 1138 FA1S $T=230020 366360 1 0 $X=230020 $Y=360940
X1930 1133 2 1128 1123 1119 1 1162 FA1S $T=234360 336120 0 0 $X=234360 $Y=335740
X1931 44 2 1138 33 40 1 59 FA1S $T=244900 366360 1 0 $X=244900 $Y=360940
X1932 1181 2 1121 1164 47 1 56 FA1S $T=249240 356280 0 0 $X=249240 $Y=355900
X1933 1212 2 55 1199 1135 1 1213 FA1S $T=259780 346200 0 0 $X=259780 $Y=345820
X1934 1215 2 1187 60 65 1 1254 FA1S $T=261020 356280 1 0 $X=261020 $Y=350860
X1935 1225 2 62 1169 1233 1 1248 FA1S $T=262880 336120 1 0 $X=262880 $Y=330700
X1936 1228 2 1118 1213 1181 1 76 FA1S $T=264120 366360 1 0 $X=264120 $Y=360940
X1937 1240 2 1151 1205 1223 1 1250 FA1S $T=267220 265560 0 0 $X=267220 $Y=265180
X1938 1241 2 1232 1230 70 1 1260 FA1S $T=267840 346200 1 0 $X=267840 $Y=340780
X1939 1245 2 1170 1236 1246 1 1264 FA1S $T=270320 285720 1 0 $X=270320 $Y=280300
X1940 1247 2 1192 1227 1226 1 1263 FA1S $T=271560 326040 0 0 $X=271560 $Y=325660
X1941 1251 2 72 1260 1212 1 1266 FA1S $T=274040 346200 0 0 $X=274040 $Y=345820
X1942 1252 2 1162 1228 1266 1 1270 FA1S $T=274660 356280 0 0 $X=274660 $Y=355900
X1943 78 2 1235 74 1190 1 1271 FA1S $T=275900 265560 1 0 $X=275900 $Y=260140
X1944 1255 2 1191 73 1243 1 1273 FA1S $T=275900 315960 0 0 $X=275900 $Y=315580
X1945 1256 2 1207 1198 1253 1 1281 FA1S $T=276520 285720 0 0 $X=276520 $Y=285340
X1946 1257 2 1203 1224 1283 1 1277 FA1S $T=276520 305880 0 0 $X=276520 $Y=305500
X1947 1258 2 1178 1167 1249 1 1268 FA1S $T=276520 315960 1 0 $X=276520 $Y=310540
X1948 1259 2 1215 1268 1225 1 1275 FA1S $T=276520 336120 1 0 $X=276520 $Y=330700
X1949 1261 2 1175 1214 1244 1 1280 FA1S $T=277760 275640 0 0 $X=277760 $Y=275260
X1950 80 2 77 1174 1231 1 1284 FA1S $T=279000 265560 0 0 $X=279000 $Y=265180
X1951 1267 2 1133 1248 1241 1 1286 FA1S $T=280240 336120 0 0 $X=280240 $Y=335740
X1952 1269 2 1254 1251 1286 1 1285 FA1S $T=281480 346200 1 0 $X=281480 $Y=340780
X1953 1272 2 1237 1220 1262 1 1293 FA1S $T=282720 295800 1 0 $X=282720 $Y=290380
X1954 1278 2 1272 1250 1245 1 1314 FA1S $T=284580 285720 1 0 $X=284580 $Y=280300
X1955 1279 2 1263 1267 1275 1 1299 FA1S $T=284580 326040 0 0 $X=284580 $Y=325660
X1956 1287 2 1247 1277 1258 1 1307 FA1S $T=287680 315960 0 0 $X=287680 $Y=315580
X1957 1288 2 85 1274 1303 1 1304 FA1S $T=288300 356280 0 0 $X=288300 $Y=355900
X1958 87 2 88 1304 82 1 84 FA1S $T=300080 366360 0 180 $X=288300 $Y=360940
X1959 1289 2 1273 1259 1307 1 1311 FA1S $T=288920 326040 1 0 $X=288920 $Y=320620
X1960 1292 2 1302 1264 1256 1 1310 FA1S $T=289540 285720 0 0 $X=289540 $Y=285340
X1961 1295 2 1255 1281 1257 1 1315 FA1S $T=290160 305880 1 0 $X=290160 $Y=300460
X1962 1296 2 1305 1287 1315 1 1319 FA1S $T=290780 305880 0 0 $X=290780 $Y=305500
X1963 1297 2 86 89 1294 1 1326 FA1S $T=291400 265560 1 0 $X=291400 $Y=260140
X1964 1294 2 1240 1284 1261 1 1317 FA1S $T=291400 265560 0 0 $X=291400 $Y=265180
X1965 1298 2 1271 1278 1317 1 1327 FA1S $T=292020 275640 1 0 $X=292020 $Y=270220
X1966 1302 2 1242 1156 1276 1 1305 FA1S $T=292640 295800 0 0 $X=292640 $Y=295420
X1967 1300 2 1282 1291 1324 1 1332 FA1S $T=293880 336120 0 0 $X=293880 $Y=335740
X1968 1308 2 1313 1300 1337 1 1321 FA1S $T=294500 336120 1 0 $X=294500 $Y=330700
X1969 1309 2 1265 1301 1334 1 1328 FA1S $T=294500 356280 1 0 $X=294500 $Y=350860
X1970 1312 2 1293 1295 1310 1 1331 FA1S $T=296360 295800 1 0 $X=296360 $Y=290380
X1971 1318 2 1280 1292 1314 1 1330 FA1S $T=298220 275640 0 0 $X=298220 $Y=275260
X1972 1325 2 1345 1332 1309 1 1353 FA1S $T=299460 346200 0 0 $X=299460 $Y=345820
X1973 1349 2 1363 1328 1288 1 90 FA1S $T=314340 356280 1 180 $X=302560 $Y=355900
X1974 1355 2 1329 1366 1348 1 1382 FA1S $T=306900 326040 1 0 $X=306900 $Y=320620
X1975 1366 2 1290 1376 1368 1 1337 FA1S $T=318680 326040 1 180 $X=306900 $Y=325660
X1976 1356 2 1379 1320 1339 1 1392 FA1S $T=307520 305880 0 0 $X=307520 $Y=305500
X1977 1371 2 1386 1444 1340 1 1344 FA1S $T=320540 295800 1 180 $X=308760 $Y=295420
X1978 1362 2 1338 1356 1344 1 1396 FA1S $T=308760 305880 1 0 $X=308760 $Y=300460
X1979 1373 2 1388 1383 1323 1 1347 FA1S $T=321160 285720 0 180 $X=309380 $Y=280300
X1980 1365 2 1342 1347 1371 1 1391 FA1S $T=309380 295800 1 0 $X=309380 $Y=290380
X1981 1374 2 1393 1343 1381 1 1348 FA1S $T=321160 315960 1 180 $X=309380 $Y=315580
X1982 1370 2 1354 1390 1373 1 1402 FA1S $T=311240 275640 0 0 $X=311240 $Y=275260
X1983 101 2 1416 1398 1359 1 1358 FA1S $T=324260 265560 0 180 $X=312480 $Y=260140
X1984 1378 2 1341 1358 1399 1 1407 FA1S $T=312480 275640 1 0 $X=312480 $Y=270220
X1985 1404 2 1441 1374 1392 1 1395 FA1S $T=321160 315960 1 0 $X=321160 $Y=310540
X1986 1399 2 1446 1449 1336 1 1390 FA1S $T=333560 285720 0 180 $X=321780 $Y=280300
X1987 1437 2 1544 1549 1540 1 1369 FA1S $T=363320 346200 1 180 $X=351540 $Y=345820
X1988 1380 2 1532 1528 1547 1 1463 FA1S $T=366420 336120 1 180 $X=354640 $Y=335740
X1989 1546 2 1559 1564 1548 1 1528 FA1S $T=367660 326040 1 180 $X=355880 $Y=325660
X1990 1474 2 1550 1563 1546 1 1475 FA1S $T=368900 326040 0 180 $X=357120 $Y=320620
X1991 1518 2 1561 1565 1553 1 1503 FA1S $T=369520 285720 0 180 $X=357740 $Y=280300
X1992 1550 2 1566 1573 1555 1 1532 FA1S $T=369520 315960 1 180 $X=357740 $Y=315580
X1993 1508 2 1574 1554 1557 1 1523 FA1S $T=370760 315960 0 180 $X=358980 $Y=310540
X1994 1530 2 1620 1545 1562 1 1511 FA1S $T=372620 305880 1 180 $X=360840 $Y=305500
X1995 1375 2 1585 1567 1556 1 1413 FA1S $T=373240 346200 0 180 $X=361460 $Y=340780
X1996 1538 2 1584 1588 1568 1 1497 FA1S $T=375100 265560 1 180 $X=363320 $Y=265180
X1997 1567 2 1578 1569 1576 1 1540 FA1S $T=376340 346200 1 180 $X=364560 $Y=345820
X1998 1569 2 1622 1611 1577 1 1551 FA1S $T=376340 356280 0 180 $X=364560 $Y=350860
X1999 1549 2 147 1551 1580 1 149 FA1S $T=364560 356280 0 0 $X=364560 $Y=355900
X2000 1565 2 1586 1593 1579 1 1545 FA1S $T=376960 285720 1 180 $X=365180 $Y=285340
X2001 146 2 1592 148 1581 1 1531 FA1S $T=377580 265560 0 180 $X=365800 $Y=260140
X2002 1562 2 1560 1596 1582 1 1554 FA1S $T=377580 295800 1 180 $X=365800 $Y=295420
X2003 1547 2 1591 1599 1558 1 1556 FA1S $T=378820 336120 0 180 $X=367040 $Y=330700
X2004 1586 2 1512 1594 1589 1 1560 FA1S $T=381300 295800 0 180 $X=369520 $Y=290380
X2005 1548 2 1602 1572 1587 1 1558 FA1S $T=382540 326040 1 180 $X=370760 $Y=325660
X2006 1590 2 1613 1605 1597 1 1571 FA1S $T=383780 275640 0 180 $X=372000 $Y=270220
X2007 1566 2 1609 1614 1598 1 1572 FA1S $T=383780 326040 0 180 $X=372000 $Y=320620
X2008 1514 2 1571 1603 1601 1 1491 FA1S $T=384400 285720 0 180 $X=372620 $Y=280300
X2009 1557 2 1617 1618 1575 1 1563 FA1S $T=384400 315960 1 180 $X=372620 $Y=315580
X2010 1574 2 1606 1604 1595 1 1575 FA1S $T=385640 315960 0 180 $X=373860 $Y=310540
X2011 1602 2 1627 1635 1610 1 1583 FA1S $T=386880 336120 1 180 $X=375100 $Y=335740
X2012 1604 2 1527 1642 1608 1 1573 FA1S $T=387500 305880 0 180 $X=375720 $Y=300460
X2013 1581 2 1631 1616 1590 1 1588 FA1S $T=388740 265560 1 180 $X=376960 $Y=265180
X2014 1585 2 1644 1583 1615 1 1544 FA1S $T=389360 346200 0 180 $X=377580 $Y=340780
X2015 1611 2 1630 1636 1621 1 150 FA1S $T=389360 356280 1 180 $X=377580 $Y=355900
X2016 1576 2 1600 1623 152 1 1580 FA1S $T=389360 366360 0 180 $X=377580 $Y=360940
X2017 1615 2 1639 1646 151 1 1577 FA1S $T=389980 346200 1 180 $X=378200 $Y=345820
X2018 1561 2 1640 1633 1612 1 1579 FA1S $T=390600 285720 1 180 $X=378820 $Y=285340
X2019 1612 2 1641 1634 1625 1 1596 FA1S $T=391220 295800 1 180 $X=379440 $Y=295420
X2020 1592 2 159 1648 158 1 1584 FA1S $T=392460 265560 0 180 $X=380680 $Y=260140
X2021 1606 2 1629 1654 1638 1 1559 FA1S $T=392460 336120 0 180 $X=380680 $Y=330700
X2022 1618 2 1664 1665 1658 1 1555 FA1S $T=399280 315960 1 180 $X=387500 $Y=315580
X2023 1662 2 1669 1670 1667 1 1617 FA1S $T=401140 315960 0 180 $X=389360 $Y=310540
X2024 1568 2 1679 1682 1671 1 1603 FA1S $T=402380 265560 1 180 $X=390600 $Y=265180
X2025 1671 2 182 1651 1656 1 1693 FA1S $T=394940 275640 1 0 $X=394940 $Y=270220
X2026 1672 2 1673 1666 1663 1 1600 FA1S $T=394940 346200 1 0 $X=394940 $Y=340780
X2027 1622 2 1680 1703 1692 1 172 FA1S $T=410440 356280 1 180 $X=398660 $Y=355900
X2028 1688 2 1699 1674 1675 1 1595 FA1S $T=400520 305880 1 0 $X=400520 $Y=300460
X2029 1658 2 1661 1686 1685 1 1587 FA1S $T=402380 315960 0 0 $X=402380 $Y=315580
X2030 1700 2 1687 1683 1698 1 1593 FA1S $T=404240 285720 1 0 $X=404240 $Y=280300
X2031 1620 2 1681 1662 1688 1 1582 FA1S $T=405480 315960 1 0 $X=405480 $Y=310540
X2032 1701 2 185 1707 1690 1 1644 FA1S $T=406720 346200 0 0 $X=406720 $Y=345820
X2033 1682 2 1705 1684 1702 1 1726 FA1S $T=407340 275640 1 0 $X=407340 $Y=270220
X2034 1564 2 1676 1701 1708 1 1591 FA1S $T=407340 336120 1 0 $X=407340 $Y=330700
X2035 1601 2 1700 1693 1726 1 1553 FA1S $T=407960 275640 0 0 $X=407960 $Y=275260
X2036 1708 2 1695 1689 1678 1 1716 FA1S $T=407960 326040 1 0 $X=407960 $Y=320620
X2037 1599 2 1709 1672 1716 1 1578 FA1S $T=419740 336120 1 180 $X=407960 $Y=335740
X2038 1709 2 1696 187 1706 1 1623 FA1S $T=408580 366360 1 0 $X=408580 $Y=360940
X2039 1718 2 1712 1728 1714 1 1743 FA1S $T=412300 285720 0 0 $X=412300 $Y=285340
X2040 1747 2 1733 1762 1718 1 1776 FA1S $T=424080 285720 1 0 $X=424080 $Y=280300
X2041 1760 2 1711 1774 1755 1 1781 FA1S $T=427800 295800 1 0 $X=427800 $Y=290380
X2042 1755 2 1753 1737 1757 1 1786 FA1S $T=428420 315960 0 0 $X=428420 $Y=315580
X2043 1769 2 1756 1746 1759 1 1788 FA1S $T=430280 336120 0 0 $X=430280 $Y=335740
X2044 1770 2 1773 1744 213 1 1802 FA1S $T=430280 356280 0 0 $X=430280 $Y=355900
X2045 1778 2 1758 1764 1769 1 1791 FA1S $T=432140 326040 1 0 $X=432140 $Y=320620
X2046 225 2 1761 1750 1787 1 1798 FA1S $T=435860 265560 0 0 $X=435860 $Y=265180
X2047 1783 2 1768 1743 1812 1 1815 FA1S $T=436480 285720 0 0 $X=436480 $Y=285340
X2048 1789 2 1775 1800 1770 1 1828 FA1S $T=438340 346200 1 0 $X=438340 $Y=340780
X2049 1790 2 1803 1781 1792 1 1811 FA1S $T=438960 305880 1 0 $X=438960 $Y=300460
X2050 1792 2 1780 1786 1807 1 1813 FA1S $T=439580 305880 0 0 $X=439580 $Y=305500
X2051 1809 2 1810 1776 1783 1 1831 FA1S $T=445780 275640 1 0 $X=445780 $Y=270220
X2052 1819 2 1794 1788 1821 1 1837 FA1S $T=448880 336120 0 0 $X=448880 $Y=335740
X2053 1822 2 1747 1798 1845 1 1852 FA1S $T=450120 265560 0 0 $X=450120 $Y=265180
X2054 1824 2 1795 1802 1847 1 1851 FA1S $T=450740 356280 0 0 $X=450740 $Y=355900
X2055 1827 2 1817 1791 1819 1 1850 FA1S $T=451360 326040 0 0 $X=451360 $Y=325660
X2056 1839 2 1830 1828 1824 1 1866 FA1S $T=455700 356280 1 0 $X=455700 $Y=350860
X2057 1858 2 1844 1871 1850 1 1832 FA1S $T=468720 326040 0 180 $X=456940 $Y=320620
X2058 1849 2 1778 1813 1843 1 1876 FA1S $T=457560 305880 0 0 $X=457560 $Y=305500
X2059 1855 2 1789 1837 1859 1 1891 FA1S $T=458180 346200 1 0 $X=458180 $Y=340780
X2060 1865 2 247 1851 1880 1 255 FA1S $T=463760 356280 0 0 $X=463760 $Y=355900
X2061 1878 2 1760 1815 1848 1 1911 FA1S $T=468100 295800 1 0 $X=468100 $Y=290380
X2062 1899 2 1856 1881 1811 1 1915 FA1S $T=474300 295800 0 0 $X=474300 $Y=295420
X2063 1903 2 1872 1898 1866 1 1918 FA1S $T=475540 356280 1 0 $X=475540 $Y=350860
X2064 1913 2 1904 1865 1918 1 1896 FA1S $T=488560 356280 1 180 $X=476780 $Y=355900
X2065 1907 2 1884 1790 1934 1 1931 FA1S $T=477400 285720 0 0 $X=477400 $Y=285340
X2066 1910 2 1892 1809 1927 1 1939 FA1S $T=479880 275640 0 0 $X=479880 $Y=275260
X2067 1919 2 1885 1827 1923 1 1942 FA1S $T=481740 315960 0 0 $X=481740 $Y=315580
X2068 1922 2 1908 1839 1938 1 1948 FA1S $T=482360 346200 1 0 $X=482360 $Y=340780
X2069 1929 2 1832 1922 1917 1 1949 FA1S $T=484220 336120 0 0 $X=484220 $Y=335740
X2070 1943 2 1855 1928 1950 1 1917 FA1S $T=498480 336120 0 180 $X=486700 $Y=330700
X2071 1940 2 1876 1858 1960 1 1958 FA1S $T=488560 326040 1 0 $X=488560 $Y=320620
X2072 1944 2 1891 1903 1948 1 1933 FA1S $T=489180 346200 0 0 $X=489180 $Y=345820
X2073 1952 2 1942 1943 1958 1 1965 FA1S $T=492900 326040 0 0 $X=492900 $Y=325660
X2074 283 2 1822 1966 1975 1 1935 FA1S $T=507160 265560 1 180 $X=495380 $Y=265180
X2075 1961 2 1849 1945 1979 1 1983 FA1S $T=495380 305880 0 0 $X=495380 $Y=305500
X2076 1963 2 1915 1919 1983 1 1984 FA1S $T=496620 315960 1 0 $X=496620 $Y=310540
X2077 1968 2 1878 1937 1993 1 1986 FA1S $T=497860 285720 1 0 $X=497860 $Y=280300
X2078 1971 2 1911 1899 1994 1 1991 FA1S $T=499100 295800 0 0 $X=499100 $Y=295420
X2079 1982 2 1852 1900 2008 1 2014 FA1S $T=502200 275640 0 0 $X=502200 $Y=275260
X2080 2001 2 2027 1931 1961 1 2032 FA1S $T=507780 305880 0 0 $X=507780 $Y=305500
X2081 2011 2 1991 1963 2032 1 2028 FA1S $T=509640 315960 1 0 $X=509640 $Y=310540
X2082 2037 2 2053 2014 1947 1 2058 FA1S $T=515840 295800 1 0 $X=515840 $Y=290380
X2083 2064 2 2050 2086 2058 1 2072 FA1S $T=523900 305880 1 0 $X=523900 $Y=300460
X2084 2085 2 2127 1939 1968 1 2050 FA1S $T=537540 285720 1 180 $X=525760 $Y=285340
X2085 2110 2 2122 1946 2085 1 2077 FA1S $T=543740 275640 0 180 $X=531960 $Y=270220
X2086 377 2 368 2258 2291 1 392 FA1S $T=577220 366360 1 0 $X=577220 $Y=360940
X2087 394 2 398 2351 403 1 395 FA1S $T=602640 366360 0 180 $X=590860 $Y=360940
X2088 2369 2 2349 2371 2438 1 2393 FA1S $T=603260 295800 0 0 $X=603260 $Y=295420
X2089 2388 2 2343 2287 2397 1 410 FA1S $T=618140 275640 0 180 $X=606360 $Y=270220
X2090 2389 2 419 2388 2393 1 411 FA1S $T=619380 265560 0 180 $X=607600 $Y=260140
X2091 2423 2 2443 2369 2429 1 2399 FA1S $T=628060 295800 0 180 $X=616280 $Y=290380
X2092 2409 2 2423 2408 2435 1 2403 FA1S $T=628680 305880 0 180 $X=616900 $Y=300460
X2093 2411 2 2211 2396 2414 1 2443 FA1S $T=616900 315960 0 0 $X=616900 $Y=315580
X2094 2387 2 2413 2416 2424 1 2391 FA1S $T=630540 275640 1 180 $X=618760 $Y=275260
X2095 2380 2 2436 2451 2442 1 2386 FA1S $T=630540 285720 1 180 $X=618760 $Y=285340
X2096 2418 2 2439 2411 2421 1 2408 FA1S $T=618760 305880 0 0 $X=618760 $Y=305500
X2097 2436 2 2448 2276 2444 1 2413 FA1S $T=631780 265560 1 180 $X=620000 $Y=265180
X2098 2455 2 2446 2469 2461 1 2439 FA1S $T=638600 315960 0 180 $X=626820 $Y=310540
X2099 2466 2 2325 2479 2475 1 2429 FA1S $T=641080 295800 1 180 $X=629300 $Y=295420
X2100 2471 2 2488 2466 2476 1 2435 FA1S $T=642320 305880 0 180 $X=630540 $Y=300460
X2101 2472 2 2316 2422 2490 1 2476 FA1S $T=633020 305880 0 0 $X=633020 $Y=305500
X2102 449 2 2459 2293 2484 1 2527 FA1S $T=644180 356280 1 0 $X=644180 $Y=350860
X2103 2488 2 2513 2524 2518 1 2442 FA1S $T=656580 285720 1 180 $X=644800 $Y=285340
X2104 2451 2 465 2523 2540 1 2424 FA1S $T=665260 265560 1 180 $X=653480 $Y=265180
X2105 2539 2 2521 2486 2504 1 2560 FA1S $T=657820 346200 0 0 $X=657820 $Y=345820
X2106 2541 2 2534 2516 2532 1 2563 FA1S $T=659060 326040 1 0 $X=659060 $Y=320620
X2107 2545 2 2560 2528 2541 1 2566 FA1S $T=659680 336120 1 0 $X=659680 $Y=330700
X2108 2555 2 2554 2512 2562 1 2421 FA1S $T=672080 295800 0 180 $X=660300 $Y=290380
X2109 2552 2 2498 2455 2555 1 2564 FA1S $T=662160 295800 0 0 $X=662160 $Y=295420
X2110 2571 2 2472 2563 2573 1 2557 FA1S $T=680140 305880 1 180 $X=668360 $Y=305500
X2111 2568 2 2506 2565 2517 1 2582 FA1S $T=668980 326040 0 0 $X=668980 $Y=325660
X2112 2574 2 2550 2539 2537 1 2589 FA1S $T=672080 346200 1 0 $X=672080 $Y=340780
X2113 2575 2 2508 2527 2569 1 2583 FA1S $T=672080 366360 1 0 $X=672080 $Y=360940
X2114 2595 2 2494 2477 2558 1 2606 FA1S $T=681380 315960 0 0 $X=681380 $Y=315580
X2115 2598 2 2582 2593 2566 1 2608 FA1S $T=683860 326040 0 0 $X=683860 $Y=325660
X2116 2607 2 2581 2585 2595 1 2593 FA1S $T=696260 326040 0 180 $X=684480 $Y=320620
X2117 2612 2 2568 2589 2607 1 2596 FA1S $T=691920 336120 1 0 $X=691920 $Y=330700
X2118 2726 2 533 2790 2775 1 2748 FA1S $T=750200 265560 1 180 $X=738420 $Y=265180
X2119 2771 2 537 544 534 1 2750 FA1S $T=750820 275640 0 180 $X=739040 $Y=270220
X2120 2768 2 2750 2748 2797 1 2792 FA1S $T=740280 275640 0 0 $X=740280 $Y=275260
X2121 549 2 550 560 555 1 2788 FA1S $T=761980 265560 0 180 $X=750200 $Y=260140
X2122 2775 2 2788 563 2815 1 2796 FA1S $T=765080 265560 1 180 $X=753300 $Y=265180
X2123 2797 2 551 2796 2822 1 2829 FA1S $T=753920 275640 0 0 $X=753920 $Y=275260
X2124 2801 2 2792 2827 2830 1 2808 FA1S $T=768180 295800 0 180 $X=756400 $Y=290380
X2125 2790 2 561 565 2842 1 2819 FA1S $T=771900 275640 0 180 $X=760120 $Y=270220
X2126 2827 2 2829 2819 2850 1 2856 FA1S $T=760740 285720 0 0 $X=760740 $Y=285340
X2127 2842 2 572 571 2852 1 2826 FA1S $T=776240 265560 0 180 $X=764460 $Y=260140
X2128 2822 2 567 2865 574 1 2836 FA1S $T=779960 265560 1 180 $X=768180 $Y=265180
X2129 2850 2 2826 566 2866 1 2867 FA1S $T=768180 275640 0 0 $X=768180 $Y=275260
X2130 2830 2 2870 2856 2873 1 2851 FA1S $T=785540 295800 0 180 $X=773760 $Y=290380
X2131 2870 2 2836 2867 584 1 2894 FA1S $T=775620 285720 1 0 $X=775620 $Y=280300
X2132 2815 2 2908 586 583 1 2865 FA1S $T=791120 265560 0 180 $X=779340 $Y=260140
X2133 2873 2 2916 2894 2895 1 2934 FA1S $T=788640 285720 0 0 $X=788640 $Y=285340
X2134 2866 2 2923 2905 598 1 2929 FA1S $T=789880 275640 0 0 $X=789880 $Y=275260
X2135 2916 2 601 2929 2922 1 2901 FA1S $T=801660 285720 0 180 $X=789880 $Y=280300
X2136 2852 2 2931 591 2930 1 2905 FA1S $T=804140 265560 1 180 $X=792360 $Y=265180
X2137 2922 2 611 2970 2955 1 2937 FA1S $T=815920 275640 0 180 $X=804140 $Y=270220
X2138 2906 2 2937 607 613 1 2945 FA1S $T=804140 275640 0 0 $X=804140 $Y=275260
X2139 2923 2 2947 631 2959 1 2970 FA1S $T=819020 275640 0 0 $X=819020 $Y=275260
X2140 2955 2 646 657 3011 1 3006 FA1S $T=825220 275640 1 0 $X=825220 $Y=270220
X2141 2946 2 666 3006 662 1 3019 FA1S $T=834520 275640 0 0 $X=834520 $Y=275260
X2142 3011 2 3016 3012 672 1 686 FA1S $T=839480 265560 1 0 $X=839480 $Y=260140
X2143 3034 2 691 3028 3052 1 3059 FA1S $T=849400 275640 1 0 $X=849400 $Y=270220
X2144 698 2 3055 3026 701 1 3028 FA1S $T=863040 265560 1 180 $X=851260 $Y=265180
X2145 3052 2 709 3065 706 1 3033 FA1S $T=865520 265560 0 180 $X=853740 $Y=260140
X2146 3032 2 3034 695 3079 1 3080 FA1S $T=856840 285720 1 0 $X=856840 $Y=280300
X2147 3079 2 3084 3059 3086 1 3057 FA1S $T=876680 275640 0 180 $X=864900 $Y=270220
X2148 3084 2 719 3033 712 1 3104 FA1S $T=868000 265560 1 0 $X=868000 $Y=260140
X2149 3086 2 731 3104 3121 1 3124 FA1S $T=879780 275640 1 0 $X=879780 $Y=270220
X2150 3121 2 3136 735 733 1 3109 FA1S $T=895280 265560 1 180 $X=883500 $Y=265180
X2151 3152 2 3155 3159 3157 1 3138 FA1S $T=909540 326040 1 180 $X=897760 $Y=325660
X2152 3157 2 3144 3205 3193 1 3087 FA1S $T=923800 326040 0 180 $X=912020 $Y=320620
X2153 3191 2 3181 3200 3190 1 3093 FA1S $T=925660 305880 0 180 $X=913880 $Y=300460
X2154 3193 2 3171 3210 3196 1 3178 FA1S $T=925660 315960 1 180 $X=913880 $Y=315580
X2155 3190 2 3175 3208 761 1 3154 FA1S $T=926280 275640 1 180 $X=914500 $Y=275260
X2156 3196 2 3164 3204 3191 1 3118 FA1S $T=926280 305880 1 180 $X=914500 $Y=305500
X2157 3279 2 3288 3270 3282 1 812 FA1S $T=964100 275640 0 180 $X=952320 $Y=270220
X2158 3278 2 3293 3295 3284 1 3268 FA1S $T=964720 295800 1 180 $X=952940 $Y=295420
X2159 3283 2 3294 3300 3289 1 817 FA1S $T=965960 265560 1 180 $X=954180 $Y=265180
X2160 3274 2 3279 3268 823 1 3213 FA1S $T=954180 285720 1 0 $X=954180 $Y=280300
X2161 3285 2 3278 3276 3274 1 3261 FA1S $T=965960 305880 0 180 $X=954180 $Y=300460
X2162 3284 2 3303 3308 3283 1 3270 FA1S $T=966580 285720 1 180 $X=954800 $Y=285340
X2163 3297 2 3312 3310 3302 1 3276 FA1S $T=970300 305880 1 180 $X=958520 $Y=305500
X2164 3282 2 3326 3341 838 1 833 FA1S $T=977740 265560 1 180 $X=965960 $Y=265180
X2165 3318 2 3297 3344 3285 1 3304 FA1S $T=978980 315960 1 180 $X=967200 $Y=315580
X2166 3321 2 3311 3330 3299 1 3308 FA1S $T=980220 285720 1 180 $X=968440 $Y=285340
X2167 3310 2 3305 3340 3324 1 3293 FA1S $T=980220 305880 0 180 $X=968440 $Y=300460
X2168 3325 2 3343 3338 3318 1 3296 FA1S $T=981460 326040 0 180 $X=969680 $Y=320620
X2169 3327 2 3345 3337 3321 1 3295 FA1S $T=982080 295800 0 180 $X=970300 $Y=290380
X2170 3347 2 3363 3352 3327 1 3312 FA1S $T=988280 315960 0 180 $X=976500 $Y=310540
X2171 3329 2 3373 3378 3358 1 3326 FA1S $T=992000 265560 1 180 $X=980220 $Y=265180
X2172 3343 2 3371 3397 3347 1 3344 FA1S $T=992620 315960 1 180 $X=980840 $Y=315580
X2173 3364 2 3381 3385 3360 1 3352 FA1S $T=994480 305880 0 180 $X=982700 $Y=300460
X2174 3360 2 3386 3393 3374 1 3345 FA1S $T=995720 295800 0 180 $X=983940 $Y=290380
X2175 3367 2 3387 3382 3379 1 3338 FA1S $T=995720 326040 1 180 $X=983940 $Y=325660
X2176 3372 2 3367 3407 3325 1 3348 FA1S $T=996340 336120 0 180 $X=984560 $Y=330700
X2177 879 2 3399 3401 3380 1 862 FA1S $T=996960 265560 0 180 $X=985180 $Y=260140
X2178 3370 2 3391 3390 3331 1 3302 FA1S $T=996960 295800 1 180 $X=985180 $Y=295420
X2179 3405 2 3418 3414 3372 1 3332 FA1S $T=1004400 336120 1 180 $X=992620 $Y=335740
X2180 3417 2 3403 3437 3364 1 3397 FA1S $T=1008740 315960 1 180 $X=996960 $Y=315580
X2181 3406 2 3422 3404 3428 1 3394 FA1S $T=1009360 295800 0 180 $X=997580 $Y=290380
X2182 3423 2 3452 3406 3417 1 3387 FA1S $T=1009980 326040 1 180 $X=998200 $Y=325660
X2183 3414 2 3444 3447 3423 1 3407 FA1S $T=1011840 336120 0 180 $X=1000060 $Y=330700
X2184 3465 2 3443 3446 3473 1 3457 FA1S $T=1014320 285720 1 0 $X=1014320 $Y=280300
X2185 3474 2 3471 3487 3465 1 3447 FA1S $T=1026100 326040 1 180 $X=1014320 $Y=325660
X2186 3479 2 3477 3468 3451 1 3493 FA1S $T=1020520 295800 1 0 $X=1020520 $Y=290380
X2187 3501 2 3503 3490 3478 1 3487 FA1S $T=1027960 326040 1 0 $X=1027960 $Y=320620
X2188 3525 2 3516 3527 3474 1 3418 FA1S $T=1038500 326040 0 0 $X=1038500 $Y=325660
X2189 1072 13 1095 2 1 XNR2HS $T=221960 326040 0 0 $X=221960 $Y=325660
X2190 7 14 15 2 1 XNR2HS $T=221960 366360 1 0 $X=221960 $Y=360940
X2191 7 25 1110 2 1 XNR2HS $T=238700 356280 1 180 $X=233120 $Y=355900
X2192 7 29 1113 2 1 XNR2HS $T=241180 356280 0 180 $X=235600 $Y=350860
X2193 21 29 1125 2 1 XNR2HS $T=242420 275640 0 180 $X=236840 $Y=270220
X2194 1140 1136 1115 2 1 XNR2HS $T=243040 315960 1 180 $X=237460 $Y=315580
X2195 1140 31 1124 2 1 XNR2HS $T=243040 336120 0 180 $X=237460 $Y=330700
X2196 1114 1136 1143 2 1 XNR2HS $T=238700 285720 0 0 $X=238700 $Y=285340
X2197 1114 1134 1147 2 1 XNR2HS $T=239320 285720 1 0 $X=239320 $Y=280300
X2198 1114 1137 1148 2 1 XNR2HS $T=239940 295800 1 0 $X=239940 $Y=290380
X2199 1117 1134 1127 2 1 XNR2HS $T=239940 315960 1 0 $X=239940 $Y=310540
X2200 34 36 1141 2 1 XNR2HS $T=246760 265560 0 180 $X=241180 $Y=260140
X2201 1155 38 1144 2 1 XNR2HS $T=246760 305880 0 180 $X=241180 $Y=300460
X2202 1155 41 1150 2 1 XNR2HS $T=248620 305880 1 180 $X=243040 $Y=305500
X2203 1140 36 1160 2 1 XNR2HS $T=243040 326040 1 0 $X=243040 $Y=320620
X2204 34 42 46 2 1 XNR2HS $T=247380 265560 1 0 $X=247380 $Y=260140
X2205 1114 1154 1176 2 1 XNR2HS $T=248000 285720 0 0 $X=248000 $Y=285340
X2206 1140 29 1177 2 1 XNR2HS $T=248620 336120 1 0 $X=248620 $Y=330700
X2207 1149 36 1131 2 1 XNR2HS $T=249240 346200 1 0 $X=249240 $Y=340780
X2208 1140 42 1182 2 1 XNR2HS $T=250480 315960 0 0 $X=250480 $Y=315580
X2209 1149 41 1183 2 1 XNR2HS $T=250480 336120 0 0 $X=250480 $Y=335740
X2210 1129 36 1184 2 1 XNR2HS $T=251100 295800 0 0 $X=251100 $Y=295420
X2211 49 1137 1180 2 1 XNR2HS $T=257920 285720 0 180 $X=252340 $Y=280300
X2212 49 1136 1188 2 1 XNR2HS $T=252960 275640 1 0 $X=252960 $Y=270220
X2213 49 1134 51 2 1 XNR2HS $T=253580 265560 1 0 $X=253580 $Y=260140
X2214 1129 38 1193 2 1 XNR2HS $T=253580 285720 0 0 $X=253580 $Y=285340
X2215 1129 42 1194 2 1 XNR2HS $T=253580 295800 1 0 $X=253580 $Y=290380
X2216 1149 38 1197 2 1 XNR2HS $T=254820 336120 1 0 $X=254820 $Y=330700
X2217 1149 42 1189 2 1 XNR2HS $T=255440 346200 1 0 $X=255440 $Y=340780
X2218 1129 1137 1200 2 1 XNR2HS $T=257300 295800 0 0 $X=257300 $Y=295420
X2219 1196 1134 1201 2 1 XNR2HS $T=257300 305880 0 0 $X=257300 $Y=305500
X2220 1196 1136 1202 2 1 XNR2HS $T=257920 315960 1 0 $X=257920 $Y=310540
X2221 49 1154 1204 2 1 XNR2HS $T=258540 285720 1 0 $X=258540 $Y=280300
X2222 1129 41 1206 2 1 XNR2HS $T=259160 285720 0 0 $X=259160 $Y=285340
X2223 1196 29 1219 2 1 XNR2HS $T=262880 305880 0 0 $X=262880 $Y=305500
X2224 1196 1159 1234 2 1 XNR2HS $T=270320 315960 0 0 $X=270320 $Y=315580
X2225 67 1195 1249 2 1 XNR2HS $T=274040 336120 0 0 $X=274040 $Y=335740
X2226 1218 1186 1253 2 1 XNR2HS $T=276520 295800 1 0 $X=276520 $Y=290380
X2227 1357 98 1372 2 1 XNR2HS $T=312480 366360 1 0 $X=312480 $Y=360940
X2228 1351 1367 1389 2 1 XNR2HS $T=316820 346200 1 0 $X=316820 $Y=340780
X2229 1428 1427 1450 2 1 XNR2HS $T=328600 326040 1 0 $X=328600 $Y=320620
X2230 1456 1453 1471 2 1 XNR2HS $T=334180 285720 1 0 $X=334180 $Y=280300
X2231 1439 1451 1467 2 1 XNR2HS $T=334800 295800 1 0 $X=334800 $Y=290380
X2232 191 1715 1710 2 1 XNR2HS $T=417880 305880 0 180 $X=412300 $Y=300460
X2233 194 1715 1717 2 1 XNR2HS $T=420980 315960 1 180 $X=415400 $Y=315580
X2234 1734 197 1720 2 1 XNR2HS $T=422840 326040 1 180 $X=417260 $Y=325660
X2235 191 193 1732 2 1 XNR2HS $T=417880 265560 1 0 $X=417880 $Y=260140
X2236 1719 1721 1733 2 1 XNR2HS $T=417880 285720 1 0 $X=417880 $Y=280300
X2237 195 197 1736 2 1 XNR2HS $T=419740 336120 0 0 $X=419740 $Y=335740
X2238 199 200 1735 2 1 XNR2HS $T=426560 346200 1 180 $X=420980 $Y=345820
X2239 204 1715 1725 2 1 XNR2HS $T=427180 305880 1 180 $X=421600 $Y=305500
X2240 204 193 1742 2 1 XNR2HS $T=429660 275640 0 180 $X=424080 $Y=270220
X2241 208 197 1741 2 1 XNR2HS $T=430280 326040 0 180 $X=424700 $Y=320620
X2242 212 1715 1724 2 1 XNR2HS $T=430900 295800 1 180 $X=425320 $Y=295420
X2243 208 193 1751 2 1 XNR2HS $T=425940 285720 0 0 $X=425940 $Y=285340
X2244 1734 1748 1754 2 1 XNR2HS $T=427180 305880 0 0 $X=427180 $Y=305500
X2245 201 200 210 2 1 XNR2HS $T=433380 366360 0 180 $X=427800 $Y=360940
X2246 195 1748 1771 2 1 XNR2HS $T=431520 315960 1 0 $X=431520 $Y=310540
X2247 215 221 1767 2 1 XNR2HS $T=438960 265560 0 180 $X=433380 $Y=260140
X2248 215 193 1763 2 1 XNR2HS $T=434620 275640 1 0 $X=434620 $Y=270220
X2249 223 1782 1777 2 1 XNR2HS $T=440820 346200 1 180 $X=435240 $Y=345820
X2250 208 221 1785 2 1 XNR2HS $T=437720 285720 1 0 $X=437720 $Y=280300
X2251 1796 1782 1784 2 1 XNR2HS $T=446400 336120 0 180 $X=440820 $Y=330700
X2252 230 1782 233 2 1 XNR2HS $T=443300 366360 1 0 $X=443300 $Y=360940
X2253 1734 221 1799 2 1 XNR2HS $T=443920 285720 1 0 $X=443920 $Y=280300
X2254 1779 1797 1793 2 1 XNR2HS $T=449500 326040 0 180 $X=443920 $Y=320620
X2255 1796 221 1801 2 1 XNR2HS $T=444540 295800 0 0 $X=444540 $Y=295420
X2256 195 221 1804 2 1 XNR2HS $T=445160 295800 1 0 $X=445160 $Y=290380
X2257 1779 1782 1805 2 1 XNR2HS $T=447020 336120 1 0 $X=447020 $Y=330700
X2258 223 1797 1814 2 1 XNR2HS $T=447640 315960 1 0 $X=447640 $Y=310540
X2259 230 231 1818 2 1 XNR2HS $T=448880 356280 1 0 $X=448880 $Y=350860
X2260 208 235 236 2 1 XNR2HS $T=449500 265560 1 0 $X=449500 $Y=260140
X2261 234 231 1820 2 1 XNR2HS $T=450120 366360 1 0 $X=450120 $Y=360940
X2262 1796 1823 1833 2 1 XNR2HS $T=453840 285720 0 0 $X=453840 $Y=285340
X2263 1734 1823 1834 2 1 XNR2HS $T=454460 275640 0 0 $X=454460 $Y=275260
X2264 1835 1836 1826 2 1 XNR2HS $T=460040 315960 1 180 $X=454460 $Y=315580
X2265 1779 1823 1838 2 1 XNR2HS $T=456320 295800 0 0 $X=456320 $Y=295420
X2266 1808 1836 1841 2 1 XNR2HS $T=456940 336120 1 0 $X=456940 $Y=330700
X2267 241 1823 1842 2 1 XNR2HS $T=461280 275640 0 0 $X=461280 $Y=275260
X2268 246 1836 1857 2 1 XNR2HS $T=463140 336120 1 0 $X=463140 $Y=330700
X2269 1864 249 1860 2 1 XNR2HS $T=469340 275640 0 180 $X=463760 $Y=270220
X2270 1796 249 250 2 1 XNR2HS $T=465000 265560 0 0 $X=465000 $Y=265180
X2271 1808 1862 1861 2 1 XNR2HS $T=470580 315960 1 180 $X=465000 $Y=315580
X2272 1835 1862 1867 2 1 XNR2HS $T=465620 315960 1 0 $X=465620 $Y=310540
X2273 1864 1823 1840 2 1 XNR2HS $T=466860 295800 0 0 $X=466860 $Y=295420
X2274 1868 1862 1877 2 1 XNR2HS $T=468720 326040 0 0 $X=468720 $Y=325660
X2275 1886 1836 1870 2 1 XNR2HS $T=474920 336120 0 180 $X=469340 $Y=330700
X2276 1779 249 1875 2 1 XNR2HS $T=469960 275640 1 0 $X=469960 $Y=270220
X2277 1868 1836 1873 2 1 XNR2HS $T=475540 336120 1 180 $X=469960 $Y=335740
X2278 251 249 254 2 1 XNR2HS $T=470580 265560 1 0 $X=470580 $Y=260140
X2279 1868 1887 1895 2 1 XNR2HS $T=473060 305880 0 0 $X=473060 $Y=305500
X2280 246 1862 1879 2 1 XNR2HS $T=480500 315960 0 180 $X=474920 $Y=310540
X2281 1901 1862 1893 2 1 XNR2HS $T=480500 336120 0 180 $X=474920 $Y=330700
X2282 1886 1862 1882 2 1 XNR2HS $T=475540 315960 0 0 $X=475540 $Y=315580
X2283 1806 256 261 2 1 XNR2HS $T=482360 265560 0 180 $X=476780 $Y=260140
X2284 1808 1912 1905 2 1 XNR2HS $T=485460 285720 0 180 $X=479880 $Y=280300
X2285 1901 1887 1906 2 1 XNR2HS $T=486080 315960 0 180 $X=480500 $Y=310540
X2286 1886 1887 1916 2 1 XNR2HS $T=482360 305880 0 0 $X=482360 $Y=305500
X2287 1864 1912 1920 2 1 XNR2HS $T=491040 275640 0 180 $X=485460 $Y=270220
X2288 246 1887 1932 2 1 XNR2HS $T=486080 295800 0 0 $X=486080 $Y=295420
X2289 1835 1912 1930 2 1 XNR2HS $T=496620 285720 1 180 $X=491040 $Y=285340
X2290 1779 1912 276 2 1 XNR2HS $T=492280 275640 1 0 $X=492280 $Y=270220
X2291 1796 1912 277 2 1 XNR2HS $T=492900 265560 1 0 $X=492900 $Y=260140
X2292 1925 1941 1954 2 1 XNR2HS $T=494140 356280 0 0 $X=494140 $Y=355900
X2293 241 281 287 2 1 XNR2HS $T=512740 265560 0 180 $X=507160 $Y=260140
X2294 1992 1988 2004 2 1 XNR2HS $T=509020 336120 0 0 $X=509020 $Y=335740
X2295 292 2016 1997 2 1 XNR2HS $T=516460 295800 1 180 $X=510880 $Y=295420
X2296 1806 281 291 2 1 XNR2HS $T=518320 265560 0 180 $X=512740 $Y=260140
X2297 274 2016 2003 2 1 XNR2HS $T=521420 275640 1 180 $X=515840 $Y=275260
X2298 1808 2036 2015 2 1 XNR2HS $T=522040 275640 0 180 $X=516460 $Y=270220
X2299 285 2016 2009 2 1 XNR2HS $T=522040 295800 1 180 $X=516460 $Y=295420
X2300 1987 2016 2026 2 1 XNR2HS $T=523280 305880 0 180 $X=517700 $Y=300460
X2301 2022 2024 2023 2 1 XNR2HS $T=517700 336120 0 0 $X=517700 $Y=335740
X2302 1835 2036 2006 2 1 XNR2HS $T=526380 265560 1 180 $X=520800 $Y=265180
X2303 2000 2036 2042 2 1 XNR2HS $T=531340 275640 0 180 $X=525760 $Y=270220
X2304 1864 2036 2030 2 1 XNR2HS $T=531960 265560 0 180 $X=526380 $Y=260140
X2305 2062 2070 2061 2 1 XNR2HS $T=530720 326040 0 0 $X=530720 $Y=325660
X2306 2096 2107 2084 2 1 XNR2HS $T=536920 326040 0 0 $X=536920 $Y=325660
X2307 2132 2134 2137 2 1 XNR2HS $T=543120 336120 1 0 $X=543120 $Y=330700
X2308 292 2161 2123 2 1 XNR2HS $T=551800 295800 0 180 $X=546220 $Y=290380
X2309 2167 2172 2149 2 1 XNR2HS $T=550560 326040 1 0 $X=550560 $Y=320620
X2310 274 2161 2147 2 1 XNR2HS $T=558000 275640 1 180 $X=552420 $Y=275260
X2311 285 2161 2125 2 1 XNR2HS $T=558000 285720 0 180 $X=552420 $Y=280300
X2312 1987 2161 2135 2 1 XNR2HS $T=558620 295800 0 180 $X=553040 $Y=290380
X2313 1808 2187 2164 2 1 XNR2HS $T=559240 275640 0 180 $X=553660 $Y=270220
X2314 1835 2187 2179 2 1 XNR2HS $T=562340 265560 1 180 $X=556760 $Y=265180
X2315 2185 2206 2188 2 1 XNR2HS $T=562340 326040 0 180 $X=556760 $Y=320620
X2316 215 281 348 2 1 XNR2HS $T=558620 295800 1 0 $X=558620 $Y=290380
X2317 2214 2210 2168 2 1 XNR2HS $T=564820 305880 0 180 $X=559240 $Y=300460
X2318 1864 2187 2219 2 1 XNR2HS $T=560480 275640 1 0 $X=560480 $Y=270220
X2319 2000 2187 2221 2 1 XNR2HS $T=561100 275640 0 0 $X=561100 $Y=275260
X2320 279 2205 2231 2 1 XNR2HS $T=564200 315960 1 0 $X=564200 $Y=310540
X2321 2040 2205 2243 2 1 XNR2HS $T=569780 315960 1 0 $X=569780 $Y=310540
X2322 292 2251 2245 2 1 XNR2HS $T=575980 275640 0 180 $X=570400 $Y=270220
X2323 361 2257 2247 2 1 XNR2HS $T=577220 285720 0 180 $X=571640 $Y=280300
X2324 285 2251 2241 2 1 XNR2HS $T=572260 275640 0 0 $X=572260 $Y=275260
X2325 2280 2278 350 2 1 XNR2HS $T=584660 336120 1 180 $X=579080 $Y=335740
X2326 274 2251 2253 2 1 XNR2HS $T=585900 265560 0 180 $X=580320 $Y=260140
X2327 2208 2285 295 2 1 XNR2HS $T=587760 285720 0 180 $X=582180 $Y=280300
X2328 2290 2289 2218 2 1 XNR2HS $T=588380 326040 1 180 $X=582800 $Y=325660
X2329 2185 2285 2296 2 1 XNR2HS $T=585280 315960 1 0 $X=585280 $Y=310540
X2330 2302 2298 2225 2 1 XNR2HS $T=590860 315960 1 180 $X=585280 $Y=315580
X2331 2303 2299 2212 2 1 XNR2HS $T=590860 336120 0 180 $X=585280 $Y=330700
X2332 2040 2285 2307 2 1 XNR2HS $T=587140 305880 0 0 $X=587140 $Y=305500
X2333 391 2251 2263 2 1 XNR2HS $T=587760 275640 1 0 $X=587760 $Y=270220
X2334 251 2305 397 2 1 XNR2HS $T=589000 265560 0 0 $X=589000 $Y=265180
X2335 2322 2318 358 2 1 XNR2HS $T=595200 346200 0 180 $X=589620 $Y=340780
X2336 279 2285 2327 2 1 XNR2HS $T=592720 305880 0 0 $X=592720 $Y=305500
X2337 215 2285 2332 2 1 XNR2HS $T=593960 285720 0 0 $X=593960 $Y=285340
X2338 2359 2356 404 2 1 XNR2HS $T=603880 356280 1 180 $X=598300 $Y=355900
X2339 1806 2305 405 2 1 XNR2HS $T=605120 265560 1 180 $X=599540 $Y=265180
X2340 241 2305 406 2 1 XNR2HS $T=606360 265560 0 180 $X=600780 $Y=260140
X2341 2249 2382 2371 2 1 XNR2HS $T=613180 315960 1 180 $X=607600 $Y=315580
X2342 2185 417 2361 2 1 XNR2HS $T=618140 366360 0 180 $X=612560 $Y=360940
X2343 2272 2404 2412 2 1 XNR2HS $T=616280 336120 1 0 $X=616280 $Y=330700
X2344 2272 420 2420 2 1 XNR2HS $T=618140 336120 0 0 $X=618140 $Y=335740
X2345 421 417 408 2 1 XNR2HS $T=624340 366360 0 180 $X=618760 $Y=360940
X2346 2419 420 2427 2 1 XNR2HS $T=620620 346200 1 0 $X=620620 $Y=340780
X2347 2419 2404 2428 2 1 XNR2HS $T=620620 346200 0 0 $X=620620 $Y=345820
X2348 2208 2432 2340 2 1 XNR2HS $T=626820 285720 0 180 $X=621240 $Y=280300
X2349 2445 420 2431 2 1 XNR2HS $T=629300 336120 1 180 $X=623720 $Y=335740
X2350 2195 2404 2449 2 1 XNR2HS $T=626200 346200 0 0 $X=626200 $Y=345820
X2351 241 2432 2406 2 1 XNR2HS $T=626820 285720 1 0 $X=626820 $Y=280300
X2352 2195 420 2450 2 1 XNR2HS $T=626820 346200 1 0 $X=626820 $Y=340780
X2353 2208 2251 2458 2 1 XNR2HS $T=630540 275640 0 0 $X=630540 $Y=275260
X2354 391 2404 432 2 1 XNR2HS $T=632400 356280 1 0 $X=632400 $Y=350860
X2355 2445 2454 2468 2 1 XNR2HS $T=633020 336120 1 0 $X=633020 $Y=330700
X2356 2482 2481 2469 2 1 XNR2HS $T=641700 315960 1 180 $X=636120 $Y=315580
X2357 2470 2483 2286 2 1 XNR2HS $T=644180 265560 0 180 $X=638600 $Y=260140
X2358 251 2489 2480 2 1 XNR2HS $T=644180 285720 1 180 $X=638600 $Y=285340
X2359 2470 2473 438 2 1 XNR2HS $T=644180 356280 1 180 $X=638600 $Y=355900
X2360 2000 2483 2457 2 1 XNR2HS $T=644800 275640 0 180 $X=639220 $Y=270220
X2361 428 2483 2493 2 1 XNR2HS $T=639840 315960 1 0 $X=639840 $Y=310540
X2362 391 2462 2487 2 1 XNR2HS $T=640460 346200 1 0 $X=640460 $Y=340780
X2363 436 2483 2465 2 1 XNR2HS $T=646660 265560 1 180 $X=641080 $Y=265180
X2364 1806 2489 2492 2 1 XNR2HS $T=641700 285720 1 0 $X=641700 $Y=280300
X2365 427 2489 2464 2 1 XNR2HS $T=648520 295800 0 180 $X=642940 $Y=290380
X2366 2040 2495 2497 2 1 XNR2HS $T=642940 346200 0 0 $X=642940 $Y=345820
X2367 2040 445 2496 2 1 XNR2HS $T=649140 326040 1 180 $X=643560 $Y=325660
X2368 2470 443 444 2 1 XNR2HS $T=645420 265560 1 0 $X=645420 $Y=260140
X2369 2470 2462 2503 2 1 XNR2HS $T=646040 346200 1 0 $X=646040 $Y=340780
X2370 428 445 2509 2 1 XNR2HS $T=648520 315960 1 0 $X=648520 $Y=310540
X2371 251 2432 2502 2 1 XNR2HS $T=649140 275640 1 0 $X=649140 $Y=270220
X2372 456 445 2505 2 1 XNR2HS $T=657200 346200 0 180 $X=651620 $Y=340780
X2373 425 445 2522 2 1 XNR2HS $T=651620 366360 1 0 $X=651620 $Y=360940
X2374 2000 457 2520 2 1 XNR2HS $T=658440 305880 1 180 $X=652860 $Y=305500
X2375 436 457 2519 2 1 XNR2HS $T=659680 295800 1 180 $X=654100 $Y=295420
X2376 2470 457 2515 2 1 XNR2HS $T=661540 265560 0 180 $X=655960 $Y=260140
X2377 1806 445 2514 2 1 XNR2HS $T=655960 275640 0 0 $X=655960 $Y=275260
X2378 2470 458 2536 2 1 XNR2HS $T=656580 285720 0 0 $X=656580 $Y=285340
X2379 456 2511 2529 2 1 XNR2HS $T=657200 336120 0 0 $X=657200 $Y=335740
X2380 425 2511 2535 2 1 XNR2HS $T=657200 366360 1 0 $X=657200 $Y=360940
X2381 1806 443 2538 2 1 XNR2HS $T=657820 285720 1 0 $X=657820 $Y=280300
X2382 2000 458 2546 2 1 XNR2HS $T=660920 305880 0 0 $X=660920 $Y=305500
X2383 436 2543 2501 2 1 XNR2HS $T=662160 275640 0 0 $X=662160 $Y=275260
X2384 436 458 2549 2 1 XNR2HS $T=662160 315960 0 0 $X=662160 $Y=315580
X2385 391 458 2551 2 1 XNR2HS $T=662780 265560 1 0 $X=662780 $Y=260140
X2386 2208 464 2556 2 1 XNR2HS $T=672080 356280 1 180 $X=666500 $Y=355900
X2387 2000 2543 2553 2 1 XNR2HS $T=670220 275640 0 0 $X=670220 $Y=275260
X2388 427 442 2567 2 1 XNR2HS $T=670220 336120 0 0 $X=670220 $Y=335740
X2389 2208 2543 2559 2 1 XNR2HS $T=677040 285720 0 180 $X=671460 $Y=280300
X2390 2208 442 2533 2 1 XNR2HS $T=671460 315960 0 0 $X=671460 $Y=315580
X2391 427 475 2576 2 1 XNR2HS $T=673940 295800 1 0 $X=673940 $Y=290380
X2392 251 2543 2579 2 1 XNR2HS $T=676420 275640 0 0 $X=676420 $Y=275260
X2393 2768 542 2784 2 1 XNR2HS $T=745860 285720 1 0 $X=745860 $Y=280300
X2394 547 2801 2794 2 1 XNR2HS $T=756400 295800 0 180 $X=750820 $Y=290380
X2395 2784 2794 2806 2 1 XNR2HS $T=752680 285720 0 0 $X=752680 $Y=285340
X2396 2806 576 2869 2 1 XNR2HS $T=776240 275640 1 0 $X=776240 $Y=270220
X2397 2813 2893 2879 2 1 XNR2HS $T=788020 275640 0 180 $X=782440 $Y=270220
X2398 2879 2869 2890 2 1 XNR2HS $T=782440 275640 0 0 $X=782440 $Y=275260
X2399 2965 2974 2980 2 1 XNR2HS $T=820880 285720 0 0 $X=820880 $Y=285340
X2400 2980 2990 2994 2 1 XNR2HS $T=827080 285720 0 0 $X=827080 $Y=285340
X2401 2890 3008 2990 2 1 XNR2HS $T=838860 285720 1 180 $X=833280 $Y=285340
X2402 2994 2998 3007 2 1 XNR2HS $T=833280 305880 1 0 $X=833280 $Y=300460
X2403 3498 3495 3339 2 1 XNR2HS $T=1031680 336120 0 180 $X=1026100 $Y=330700
X2404 1513 112 119 1 2 1496 OA12 $T=350920 336120 0 180 $X=347200 $Y=330700
X2405 1512 138 1527 1 2 1534 OA12 $T=364560 295800 0 180 $X=360840 $Y=290380
X2406 2603 2587 2584 1 2 2578 OA12 $T=684480 275640 0 180 $X=680760 $Y=270220
X2407 2999 2976 2988 1 2 2979 OA12 $T=829560 346200 0 180 $X=825840 $Y=340780
X2408 3457 3429 3454 1 2 3452 OA12 $T=1018040 326040 0 180 $X=1014320 $Y=320620
X2409 3493 3501 3495 1 2 3516 OA12 $T=1031680 326040 0 0 $X=1031680 $Y=325660
X2410 3492 3507 3519 1 2 3527 OA12 $T=1044080 305880 1 180 $X=1040360 $Y=305500
X2411 3595 3560 3612 1 2 3613 OA12 $T=1067020 315960 0 0 $X=1067020 $Y=315580
X2412 20 1 1110 19 1104 15 2 OAI22S $T=231880 356280 1 180 $X=228160 $Y=355900
X2413 20 1 1113 19 1102 1110 2 OAI22S $T=234980 356280 0 180 $X=231260 $Y=350860
X2414 1101 1 1115 1111 1112 1095 2 OAI22S $T=235600 326040 1 180 $X=231880 $Y=325660
X2415 1101 1 1095 1109 1121 1124 2 OAI22S $T=233120 336120 1 0 $X=233120 $Y=330700
X2416 1139 1 1127 1111 1123 1115 2 OAI22S $T=239940 326040 1 180 $X=236220 $Y=325660
X2417 20 1 1131 19 1128 1113 2 OAI22S $T=240560 346200 0 180 $X=236840 $Y=340780
X2418 1132 1 1125 1120 1153 1147 2 OAI22S $T=243040 275640 1 0 $X=243040 $Y=270220
X2419 27 1 1141 1120 1151 1125 2 OAI22S $T=247380 265560 1 180 $X=243660 $Y=265180
X2420 1157 1 19 1152 37 1146 2 OAI22S $T=247380 346200 1 180 $X=243660 $Y=345820
X2421 1132 1 1147 1158 1156 1143 2 OAI22S $T=244280 285720 0 0 $X=244280 $Y=285340
X2422 1132 1 1143 1158 1165 1148 2 OAI22S $T=246140 295800 1 0 $X=246140 $Y=290380
X2423 1166 1 1111 1161 1164 1139 2 OAI22S $T=251100 326040 1 180 $X=247380 $Y=325660
X2424 48 1 1158 1168 1167 1132 2 OAI22S $T=252340 275640 0 180 $X=248620 $Y=270220
X2425 1166 1 1139 1172 1175 1150 2 OAI22S $T=248620 315960 1 0 $X=248620 $Y=310540
X2426 1171 1 1150 1172 1170 1144 2 OAI22S $T=252960 305880 1 180 $X=249240 $Y=305500
X2427 1132 1 1148 1158 1178 1176 2 OAI22S $T=249860 295800 1 0 $X=249860 $Y=290380
X2428 27 1 46 43 1174 1141 2 OAI22S $T=254200 265560 1 180 $X=250480 $Y=265180
X2429 1171 1 1177 1172 1179 1127 2 OAI22S $T=256060 326040 0 180 $X=252340 $Y=320620
X2430 1171 1 1144 1172 1186 1182 2 OAI22S $T=252960 305880 0 0 $X=252960 $Y=305500
X2431 1146 1 1189 1173 1187 1131 2 OAI22S $T=258540 346200 1 180 $X=254820 $Y=345820
X2432 1171 1 1182 1111 1191 1160 2 OAI22S $T=259780 315960 1 180 $X=256060 $Y=315580
X2433 1171 1 1160 1111 1192 1177 2 OAI22S $T=259780 326040 0 180 $X=256060 $Y=320620
X2434 1146 1 1197 1173 1195 1189 2 OAI22S $T=260400 336120 1 180 $X=256680 $Y=335740
X2435 52 1 53 1185 1198 57 2 OAI22S $T=257920 265560 0 0 $X=257920 $Y=265180
X2436 57 1 1188 53 1208 1180 2 OAI22S $T=261020 275640 1 0 $X=261020 $Y=270220
X2437 1146 1 1183 1173 1203 1197 2 OAI22S $T=264740 336120 1 180 $X=261020 $Y=335740
X2438 57 1 51 53 1205 1188 2 OAI22S $T=265360 265560 1 180 $X=261640 $Y=265180
X2439 57 1 1180 53 1207 1204 2 OAI22S $T=265980 275640 1 180 $X=262260 $Y=275260
X2440 1222 1 1202 1211 1210 1200 2 OAI22S $T=266600 315960 1 180 $X=262880 $Y=315580
X2441 1217 1 1193 1216 1214 1194 2 OAI22S $T=268460 285720 1 180 $X=264740 $Y=285340
X2442 1157 1 1146 1173 1218 1183 2 OAI22S $T=269080 336120 1 180 $X=265360 $Y=335740
X2443 1222 1 1200 1211 1232 1234 2 OAI22S $T=266600 315960 0 0 $X=266600 $Y=315580
X2444 1222 1 1201 1211 1227 1202 2 OAI22S $T=271560 315960 0 180 $X=267840 $Y=310540
X2445 1217 1 1206 1216 1231 1193 2 OAI22S $T=272180 285720 1 180 $X=268460 $Y=285340
X2446 1217 1 1194 1216 1237 1184 2 OAI22S $T=268460 295800 1 0 $X=268460 $Y=290380
X2447 1222 1 1219 1211 1238 1201 2 OAI22S $T=274040 305880 0 180 $X=270320 $Y=300460
X2448 1222 1 1184 1211 1242 1219 2 OAI22S $T=275280 295800 1 180 $X=271560 $Y=295420
X2449 58 1 66 69 1235 1221 2 OAI22S $T=275900 265560 0 180 $X=272180 $Y=260140
X2450 1229 1 1217 1216 68 1206 2 OAI22S $T=275900 285720 1 180 $X=272180 $Y=285340
X2451 1229 1 1211 1239 1230 1222 2 OAI22S $T=275900 305880 1 180 $X=272180 $Y=305500
X2452 1481 1 1489 115 1490 1502 2 OAI22S $T=344100 346200 0 0 $X=344100 $Y=345820
X2453 1516 1 1481 1526 1501 132 2 OAI22S $T=353400 356280 1 0 $X=353400 $Y=350860
X2454 1722 1 1724 1723 1721 1710 2 OAI22S $T=421600 305880 0 180 $X=417880 $Y=300460
X2455 1722 1 1710 1723 1728 1725 2 OAI22S $T=417880 305880 0 0 $X=417880 $Y=305500
X2456 1722 1 1725 1729 1727 1717 2 OAI22S $T=418500 315960 1 0 $X=418500 $Y=310540
X2457 1722 1 1717 1723 1737 1741 2 OAI22S $T=421600 315960 0 0 $X=421600 $Y=315580
X2458 196 1 1736 1729 1738 1735 2 OAI22S $T=421600 346200 1 0 $X=421600 $Y=340780
X2459 196 1 1741 1729 1739 1720 2 OAI22S $T=427180 326040 1 180 $X=423460 $Y=325660
X2460 196 1 1735 205 1744 210 2 OAI22S $T=424080 356280 0 0 $X=424080 $Y=355900
X2461 1749 1 206 203 202 1732 2 OAI22S $T=428420 265560 0 180 $X=424700 $Y=260140
X2462 196 1 1720 1729 1746 1736 2 OAI22S $T=425320 336120 0 0 $X=425320 $Y=335740
X2463 1749 1 1732 203 1761 1742 2 OAI22S $T=430280 265560 0 0 $X=430280 $Y=265180
X2464 1749 1 1742 203 1762 1763 2 OAI22S $T=430280 275640 1 0 $X=430280 $Y=270220
X2465 1749 1 1763 1766 1768 1751 2 OAI22S $T=432140 285720 0 0 $X=432140 $Y=285340
X2466 1749 1 1751 1766 1774 1754 2 OAI22S $T=433380 295800 0 0 $X=433380 $Y=295420
X2467 216 1 1754 1766 1780 1771 2 OAI22S $T=435860 305880 0 0 $X=435860 $Y=305500
X2468 216 1 1771 1766 1764 1784 2 OAI22S $T=437720 315960 1 0 $X=437720 $Y=310540
X2469 224 1 226 1767 228 229 2 OAI22S $T=439580 265560 1 0 $X=439580 $Y=260140
X2470 227 1 1767 1785 1787 229 2 OAI22S $T=440820 275640 1 0 $X=440820 $Y=270220
X2471 216 1 1784 232 1794 1805 2 OAI22S $T=443300 336120 0 0 $X=443300 $Y=335740
X2472 216 1 1777 232 1795 233 2 OAI22S $T=443300 356280 1 0 $X=443300 $Y=350860
X2473 216 1 1805 232 1800 1777 2 OAI22S $T=451360 346200 1 180 $X=447640 $Y=345820
X2474 1816 1 1785 1799 1810 229 2 OAI22S $T=453840 275640 1 180 $X=450120 $Y=275260
X2475 1816 1 1799 1804 1812 229 2 OAI22S $T=453840 285720 0 180 $X=450120 $Y=280300
X2476 227 1 1793 1814 1817 237 2 OAI22S $T=450120 326040 1 0 $X=450120 $Y=320620
X2477 1816 1 1801 1793 1807 237 2 OAI22S $T=451980 305880 0 0 $X=451980 $Y=305500
X2478 1816 1 1804 1801 1803 237 2 OAI22S $T=452600 295800 0 0 $X=452600 $Y=295420
X2479 227 1 1814 1818 1821 237 2 OAI22S $T=456940 336120 0 180 $X=453220 $Y=330700
X2480 240 1 1818 1820 1830 238 2 OAI22S $T=460040 366360 0 180 $X=456320 $Y=360940
X2481 239 1 236 1834 242 243 2 OAI22S $T=457560 265560 1 0 $X=457560 $Y=260140
X2482 1825 1 1834 1842 1845 243 2 OAI22S $T=458800 275640 1 0 $X=458800 $Y=270220
X2483 1825 1 1833 1838 1848 1854 2 OAI22S $T=459420 295800 1 0 $X=459420 $Y=290380
X2484 1825 1 1840 1826 1843 1854 2 OAI22S $T=459420 315960 1 0 $X=459420 $Y=310540
X2485 1825 1 1842 1833 1853 1854 2 OAI22S $T=460040 285720 0 0 $X=460040 $Y=285340
X2486 1829 1 1826 1841 1844 1854 2 OAI22S $T=460660 315960 0 0 $X=460660 $Y=315580
X2487 240 1 1820 244 1847 238 2 OAI22S $T=464380 366360 0 180 $X=460660 $Y=360940
X2488 1829 1 1841 1857 1859 1854 2 OAI22S $T=461280 336120 0 0 $X=461280 $Y=335740
X2489 1825 1 1838 1840 1856 1854 2 OAI22S $T=466240 295800 1 180 $X=462520 $Y=295420
X2490 1829 1 1857 1870 1872 1883 2 OAI22S $T=468100 346200 0 0 $X=468100 $Y=345820
X2491 1829 1 1870 1873 1880 1883 2 OAI22S $T=469960 356280 1 0 $X=469960 $Y=350860
X2492 1869 1 1875 1860 1874 1889 2 OAI22S $T=470580 275640 0 0 $X=470580 $Y=275260
X2493 1869 1 1860 1867 1884 1889 2 OAI22S $T=471200 285720 0 0 $X=471200 $Y=285340
X2494 1869 1 1867 1861 1881 1890 2 OAI22S $T=471200 305880 1 0 $X=471200 $Y=300460
X2495 1869 1 1861 1879 1885 1890 2 OAI22S $T=471200 315960 0 0 $X=471200 $Y=315580
X2496 1869 1 1879 1882 1871 1890 2 OAI22S $T=471200 326040 1 0 $X=471200 $Y=320620
X2497 1829 1 1873 252 253 1883 2 OAI22S $T=471200 366360 1 0 $X=471200 $Y=360940
X2498 1869 1 250 1875 1892 1889 2 OAI22S $T=478640 275640 1 180 $X=474920 $Y=275260
X2499 1894 1 1877 1893 1898 1890 2 OAI22S $T=475540 336120 0 0 $X=475540 $Y=335740
X2500 1894 1 1882 1877 1908 1890 2 OAI22S $T=479260 326040 1 0 $X=479260 $Y=320620
X2501 265 1 1890 1909 1904 268 2 OAI22S $T=479880 336120 0 0 $X=479880 $Y=335740
X2502 1921 1 1920 1924 1927 1930 2 OAI22S $T=486080 285720 1 0 $X=486080 $Y=280300
X2503 1926 1 1916 1924 1923 1895 2 OAI22S $T=489800 315960 0 180 $X=486080 $Y=310540
X2504 1921 1 1905 1924 1934 1932 2 OAI22S $T=487940 295800 1 0 $X=487940 $Y=290380
X2505 1921 1 1895 1924 1928 1906 2 OAI22S $T=493520 315960 0 180 $X=489800 $Y=310540
X2506 1921 1 1930 1924 1937 1905 2 OAI22S $T=494140 285720 0 180 $X=490420 $Y=280300
X2507 1921 1 1932 1924 1945 1916 2 OAI22S $T=491660 305880 0 0 $X=491660 $Y=305500
X2508 278 1 276 282 1966 1920 2 OAI22S $T=499100 275640 1 0 $X=499100 $Y=270220
X2509 1964 1 1997 1999 1994 2009 2 OAI22S $T=509640 305880 1 0 $X=509640 $Y=300460
X2510 2002 1 2003 1999 1993 1997 2 OAI22S $T=514600 285720 0 180 $X=510880 $Y=280300
X2511 2002 1 2006 2010 1975 2015 2 OAI22S $T=512120 265560 0 0 $X=512120 $Y=265180
X2512 2002 1 2015 2010 2008 2003 2 OAI22S $T=516460 275640 0 180 $X=512740 $Y=270220
X2513 1964 1 2009 1999 1979 2026 2 OAI22S $T=513980 305880 1 0 $X=513980 $Y=300460
X2514 2002 1 2030 2010 294 2006 2 OAI22S $T=516460 265560 0 0 $X=516460 $Y=265180
X2515 2002 1 295 2010 298 2042 2 OAI22S $T=518320 265560 1 0 $X=518320 $Y=260140
X2516 2002 1 2042 2010 302 2030 2 OAI22S $T=522040 265560 1 0 $X=522040 $Y=260140
X2517 2046 1 2123 2126 2127 2125 2 OAI22S $T=540640 285720 1 0 $X=540640 $Y=280300
X2518 2046 1 2125 2126 2102 2135 2 OAI22S $T=541260 295800 0 0 $X=541260 $Y=295420
X2519 2046 1 2147 2126 2108 2123 2 OAI22S $T=548700 285720 0 180 $X=544980 $Y=280300
X2520 2151 1 2126 2146 2093 2046 2 OAI22S $T=548700 295800 1 180 $X=544980 $Y=295420
X2521 2166 1 2164 2160 332 2147 2 OAI22S $T=551800 275640 0 180 $X=548080 $Y=270220
X2522 2166 1 2219 2160 351 2179 2 OAI22S $T=566060 265560 1 180 $X=562340 $Y=265180
X2523 2220 1 2231 2222 354 348 2 OAI22S $T=568540 305880 1 180 $X=564820 $Y=305500
X2524 2166 1 2221 2160 359 2219 2 OAI22S $T=569780 265560 1 180 $X=566060 $Y=265180
X2525 364 1 2222 2234 1950 2220 2 OAI22S $T=569780 326040 0 180 $X=566060 $Y=320620
X2526 2202 1 2241 2244 2101 2247 2 OAI22S $T=568540 275640 0 0 $X=568540 $Y=275260
X2527 2220 1 2243 2222 2238 2231 2 OAI22S $T=572260 305880 1 180 $X=568540 $Y=305500
X2528 2202 1 2245 2244 2237 2241 2 OAI22S $T=569780 265560 0 0 $X=569780 $Y=265180
X2529 2220 1 2188 2222 2249 2243 2 OAI22S $T=570400 315960 0 0 $X=570400 $Y=315580
X2530 2202 1 2253 2244 372 2245 2 OAI22S $T=575980 265560 0 180 $X=572260 $Y=260140
X2531 2202 1 2263 2244 376 2253 2 OAI22S $T=579700 265560 0 180 $X=575980 $Y=260140
X2532 381 1 2269 2261 2021 1964 2 OAI22S $T=581560 326040 0 180 $X=577840 $Y=320620
X2533 2266 1 2244 2273 2122 388 2 OAI22S $T=581560 275640 0 0 $X=581560 $Y=275260
X2534 2202 1 2286 2244 389 2263 2 OAI22S $T=585280 265560 0 0 $X=585280 $Y=265180
X2535 2270 1 2296 2313 2316 2307 2 OAI22S $T=590240 305880 1 0 $X=590240 $Y=300460
X2536 396 1 2307 2313 2325 2327 2 OAI22S $T=593340 295800 0 0 $X=593340 $Y=295420
X2537 2166 1 2340 2160 400 2221 2 OAI22S $T=600780 265560 0 180 $X=597060 $Y=260140
X2538 396 1 2332 401 2343 405 2 OAI22S $T=597060 275640 1 0 $X=597060 $Y=270220
X2539 396 1 2327 2313 2349 2332 2 OAI22S $T=597680 295800 0 0 $X=597680 $Y=295420
X2540 2361 1 409 407 2351 408 2 OAI22S $T=611320 366360 0 180 $X=607600 $Y=360940
X2541 2352 1 2406 2400 418 2340 2 OAI22S $T=620620 285720 0 180 $X=616900 $Y=280300
X2542 2420 1 2425 2426 2382 2431 2 OAI22S $T=622480 336120 1 0 $X=622480 $Y=330700
X2543 2427 1 2425 2426 2440 2420 2 OAI22S $T=629920 336120 0 180 $X=626200 $Y=330700
X2544 2450 1 2425 2426 2446 2427 2 OAI22S $T=633640 336120 1 180 $X=629920 $Y=335740
X2545 2453 1 2457 2460 430 2465 2 OAI22S $T=633020 265560 0 0 $X=633020 $Y=265180
X2546 2453 1 2458 2460 2456 2457 2 OAI22S $T=633020 275640 1 0 $X=633020 $Y=270220
X2547 2467 1 2464 2460 2438 2458 2 OAI22S $T=637980 295800 0 180 $X=634260 $Y=290380
X2548 2478 1 435 434 2448 431 2 OAI22S $T=639220 346200 1 180 $X=635500 $Y=345820
X2549 2453 1 2465 2460 437 2286 2 OAI22S $T=636740 265560 0 0 $X=636740 $Y=265180
X2550 2487 1 2425 2426 2477 2450 2 OAI22S $T=641700 336120 1 180 $X=637980 $Y=335740
X2551 2467 1 2480 2460 2475 2464 2 OAI22S $T=642320 295800 0 180 $X=638600 $Y=290380
X2552 432 1 2452 439 2484 2449 2 OAI22S $T=638600 356280 1 0 $X=638600 $Y=350860
X2553 2485 1 2452 439 2481 2474 2 OAI22S $T=642940 326040 0 180 $X=639220 $Y=320620
X2554 2449 1 2452 439 2486 2428 2 OAI22S $T=639220 346200 0 0 $X=639220 $Y=345820
X2555 2412 1 2452 439 2482 2468 2 OAI22S $T=643560 336120 0 180 $X=639840 $Y=330700
X2556 2453 1 2492 402 2490 2480 2 OAI22S $T=645420 295800 1 180 $X=641700 $Y=295420
X2557 2428 1 2452 439 2491 2412 2 OAI22S $T=646040 336120 1 180 $X=642320 $Y=335740
X2558 2467 1 2493 402 2498 2492 2 OAI22S $T=649760 305880 0 180 $X=646040 $Y=300460
X2559 2507 1 2501 378 2397 444 2 OAI22S $T=650380 265560 1 180 $X=646660 $Y=265180
X2560 2352 1 2502 2400 447 2406 2 OAI22S $T=651000 285720 0 180 $X=647280 $Y=280300
X2561 452 1 450 2500 448 446 2 OAI22S $T=651620 315960 1 180 $X=647900 $Y=315580
X2562 441 1 435 434 2508 2503 2 OAI22S $T=647900 366360 1 0 $X=647900 $Y=360940
X2563 2352 1 2505 2510 2512 2509 2 OAI22S $T=649140 305880 0 0 $X=649140 $Y=305500
X2564 2503 1 2425 434 2504 2487 2 OAI22S $T=652860 336120 1 180 $X=649140 $Y=335740
X2565 2352 1 2509 2510 2513 2514 2 OAI22S $T=649760 295800 1 0 $X=649760 $Y=290380
X2566 455 1 2515 454 2444 451 2 OAI22S $T=655340 265560 0 180 $X=651620 $Y=260140
X2567 2381 1 2496 2510 2516 2505 2 OAI22S $T=656580 326040 0 180 $X=652860 $Y=320620
X2568 2381 1 2522 2510 2517 2496 2 OAI22S $T=656580 326040 1 180 $X=652860 $Y=325660
X2569 2519 1 455 454 2524 2515 2 OAI22S $T=653480 295800 1 0 $X=653480 $Y=290380
X2570 2352 1 2514 2510 2523 2502 2 OAI22S $T=657820 285720 0 180 $X=654100 $Y=280300
X2571 455 1 2520 450 2461 2519 2 OAI22S $T=654720 315960 1 0 $X=654720 $Y=310540
X2572 2530 1 2529 402 2528 2493 2 OAI22S $T=660300 326040 1 180 $X=656580 $Y=325660
X2573 446 1 2533 450 2532 2520 2 OAI22S $T=661540 315960 1 180 $X=657820 $Y=315580
X2574 2530 1 2535 2531 459 2497 2 OAI22S $T=661540 356280 1 180 $X=657820 $Y=355900
X2575 2530 1 2497 2531 2537 2529 2 OAI22S $T=662780 356280 0 180 $X=659060 $Y=350860
X2576 2536 1 2547 466 2554 2551 2 OAI22S $T=664640 285720 0 0 $X=664640 $Y=285340
X2577 2556 1 461 467 2550 2546 2 OAI22S $T=668980 346200 0 180 $X=665260 $Y=340780
X2578 468 1 469 467 471 2556 2 OAI22S $T=666500 366360 1 0 $X=666500 $Y=360940
X2579 2507 1 2553 378 2540 2501 2 OAI22S $T=670840 275640 0 180 $X=667120 $Y=270220
X2580 2507 1 2559 470 2518 2553 2 OAI22S $T=670840 285720 0 180 $X=667120 $Y=280300
X2581 2549 1 461 467 2558 2536 2 OAI22S $T=671460 315960 1 180 $X=667740 $Y=315580
X2582 2551 1 2547 466 2479 472 2 OAI22S $T=668980 265560 1 0 $X=668980 $Y=260140
X2583 2546 1 461 467 2565 2549 2 OAI22S $T=676420 326040 0 180 $X=672700 $Y=320620
X2584 446 1 473 450 2569 2567 2 OAI22S $T=676420 356280 1 180 $X=672700 $Y=355900
X2585 2507 1 2576 470 2562 2559 2 OAI22S $T=679520 285720 1 180 $X=675800 $Y=285340
X2586 478 1 477 476 2570 2538 2 OAI22S $T=680760 356280 1 180 $X=677040 $Y=355900
X2587 446 1 2567 450 2581 2533 2 OAI22S $T=677660 326040 1 0 $X=677660 $Y=320620
X2588 2507 1 2538 378 2585 2579 2 OAI22S $T=679520 285720 0 0 $X=679520 $Y=285340
X2589 478 1 2579 470 2594 2576 2 OAI22S $T=682620 295800 1 0 $X=682620 $Y=290380
X2590 2652 1 2640 2651 2647 2617 2 OAI22S $T=708660 295800 1 180 $X=704940 $Y=295420
X2591 2682 1 512 2695 2645 2659 2 OAI22S $T=723540 336120 1 180 $X=719820 $Y=335740
X2592 2671 1 2659 2705 2661 2677 2 OAI22S $T=724160 326040 1 180 $X=720440 $Y=325660
X2593 2908 1 2921 2908 2931 2918 2 OAI22S $T=799800 265560 1 0 $X=799800 $Y=260140
X2594 2930 1 2950 2930 2947 2944 2 OAI22S $T=811580 265560 1 180 $X=807860 $Y=265180
X2595 3299 1 3301 3299 3300 3309 2 OAI22S $T=965340 275640 0 0 $X=965340 $Y=275260
X2596 3305 1 3306 3305 3311 3307 2 OAI22S $T=967200 295800 0 0 $X=967200 $Y=295420
X2597 3289 1 3314 3289 845 3316 2 OAI22S $T=969680 265560 1 0 $X=969680 $Y=260140
X2598 3294 1 3323 3294 852 3335 2 OAI22S $T=975260 265560 1 0 $X=975260 $Y=260140
X2599 3331 1 3336 3331 3340 3342 2 OAI22S $T=977740 295800 0 0 $X=977740 $Y=295420
X2600 3403 1 3408 3403 3363 3412 2 OAI22S $T=999440 315960 1 0 $X=999440 $Y=310540
X2601 3429 1 3431 3429 3437 3442 2 OAI22S $T=1006880 315960 1 0 $X=1006880 $Y=310540
X2602 3471 1 3426 3471 3379 3466 2 OAI22S $T=1022380 326040 0 180 $X=1018660 $Y=320620
X2603 3492 1 3494 3492 3490 3489 2 OAI22S $T=1031680 305880 1 180 $X=1027960 $Y=305500
X2604 3507 1 3500 3507 3503 3480 2 OAI22S $T=1035400 315960 0 180 $X=1031680 $Y=310540
X2605 949 1 3518 3523 3524 3526 2 OAI22S $T=1036640 265560 0 0 $X=1036640 $Y=265180
X2606 3526 1 3521 3523 3553 975 2 OAI22S $T=1049040 275640 1 0 $X=1049040 $Y=270220
X2607 972 1 3528 980 3555 983 2 OAI22S $T=1050280 265560 1 0 $X=1050280 $Y=260140
X2608 3597 1 3547 3559 3545 3588 2 OAI22S $T=1067020 295800 1 180 $X=1063300 $Y=295420
X2609 3616 1 3619 3607 3621 3633 2 OAI22S $T=1069500 305880 1 0 $X=1069500 $Y=300460
X2610 2708 2745 535 2 2760 539 1 AO22 $T=738420 366360 1 0 $X=738420 $Y=360940
X2611 2721 2749 2763 2 2766 539 1 AO22 $T=740900 346200 1 0 $X=740900 $Y=340780
X2612 2783 2728 2763 2 2777 2780 1 AO22 $T=748960 336120 1 0 $X=748960 $Y=330700
X2613 2787 2804 2800 2 2809 2780 1 AO22 $T=753920 346200 0 0 $X=753920 $Y=345820
X2614 2785 2786 2763 2 2812 2780 1 AO22 $T=755160 336120 1 0 $X=755160 $Y=330700
X2615 2811 2791 2800 2 2825 2780 1 AO22 $T=761360 336120 1 0 $X=761360 $Y=330700
X2616 2832 2840 2800 2 2843 2780 1 AO22 $T=766940 346200 0 0 $X=766940 $Y=345820
X2617 2824 2841 2800 2 2846 2780 1 AO22 $T=767560 336120 1 0 $X=767560 $Y=330700
X2618 1171 1172 1166 1 2 1190 AO12 $T=252960 315960 1 0 $X=252960 $Y=310540
X2619 1146 1173 1157 1 2 1220 AO12 $T=261640 346200 1 0 $X=261640 $Y=340780
X2620 1217 1216 1229 1 2 71 AO12 $T=272180 295800 1 0 $X=272180 $Y=290380
X2621 1541 1536 1526 1 2 135 AO12 $T=361460 356280 1 180 $X=357740 $Y=355900
X2622 1722 1729 1724 1 2 1740 AO12 $T=421600 305880 1 0 $X=421600 $Y=300460
X2623 1749 203 206 1 2 214 AO12 $T=429040 265560 1 0 $X=429040 $Y=260140
X2624 2220 2222 2188 1 2 2211 AO12 $T=566680 315960 1 180 $X=562960 $Y=315580
X2625 2270 2313 2296 1 2 2338 AO12 $T=594580 305880 1 0 $X=594580 $Y=300460
X2626 409 407 2361 1 2 2291 AO12 $T=606980 366360 0 180 $X=603260 $Y=360940
X2627 2381 2510 2522 1 2 2525 AO12 $T=653480 336120 0 0 $X=653480 $Y=335740
X2628 2530 2531 2535 1 2 463 AO12 $T=661540 356280 0 0 $X=661540 $Y=355900
X2629 2714 2715 2659 1 2 2688 AO12 $T=727880 326040 1 180 $X=724160 $Y=325660
X2630 3568 3617 3622 1 2 3620 AO12 $T=1068880 326040 0 0 $X=1068880 $Y=325660
X2631 3748 3741 3720 1 2 3643 AO12 $T=1106080 326040 0 180 $X=1102360 $Y=320620
X2632 3747 3756 3762 1 2 3755 AO12 $T=1112280 315960 1 180 $X=1108560 $Y=315580
X2633 91 93 2 1335 1 94 AOI12HS $T=303800 366360 1 0 $X=303800 $Y=360940
X2634 269 273 2 275 1 1951 AOI12HS $T=491660 366360 1 0 $X=491660 $Y=360940
X2635 1970 1973 2 1985 1 1981 AOI12HS $T=504680 336120 1 0 $X=504680 $Y=330700
X2636 2017 2024 2 2029 1 2044 AOI12HS $T=518320 336120 1 0 $X=518320 $Y=330700
X2637 2029 2048 2 2060 1 2063 AOI12HS $T=525760 326040 1 0 $X=525760 $Y=320620
X2638 2066 2070 2 2088 1 2097 AOI12HS $T=531960 326040 1 0 $X=531960 $Y=320620
X2639 2099 2107 2 2120 1 2124 AOI12HS $T=538160 326040 1 0 $X=538160 $Y=320620
X2640 2120 2119 2 2106 1 2116 AOI12HS $T=543120 315960 1 180 $X=538780 $Y=315580
X2641 2229 2210 2 2209 1 2194 AOI12HS $T=566060 295800 1 180 $X=561720 $Y=295420
X2642 2240 2210 2 2250 1 2255 AOI12HS $T=570400 295800 0 0 $X=570400 $Y=295420
X2643 2210 2268 2 2274 1 2277 AOI12HS $T=579080 305880 1 0 $X=579080 $Y=300460
X2644 2331 2337 2 2346 1 2300 AOI12HS $T=597060 326040 0 0 $X=597060 $Y=325660
X2645 2355 2358 2 2362 1 2328 AOI12HS $T=602020 346200 1 0 $X=602020 $Y=340780
X2646 2350 2358 2 2366 1 2324 AOI12HS $T=603260 336120 0 0 $X=603260 $Y=335740
X2647 2335 2358 2 2367 1 2353 AOI12HS $T=603260 356280 1 0 $X=603260 $Y=350860
X2648 2967 2969 2 2959 1 629 AOI12HS $T=820880 265560 1 180 $X=816540 $Y=265180
X2649 2992 3000 2 653 1 3012 AOI12HS $T=832040 265560 1 0 $X=832040 $Y=260140
X2650 3017 3015 2 3016 1 3026 AOI12HS $T=845680 265560 0 0 $X=845680 $Y=265180
X2651 3074 3069 2 3055 1 3065 AOI12HS $T=869860 265560 1 180 $X=865520 $Y=265180
X2652 31 2 1101 30 1 AN2B1S $T=242420 356280 1 180 $X=239320 $Y=355900
X2653 1159 2 1132 1169 1 AN2B1S $T=247380 295800 0 0 $X=247380 $Y=295420
X2654 1159 2 1145 1199 1 AN2B1S $T=262880 315960 1 180 $X=259780 $Y=315580
X2655 1154 2 57 1224 1 AN2B1S $T=264740 285720 1 0 $X=264740 $Y=280300
X2656 1159 2 66 1236 1 AN2B1S $T=267220 275640 0 0 $X=267220 $Y=275260
X2657 1252 2 83 1282 1 AN2B1S $T=287060 356280 1 0 $X=287060 $Y=350860
X2658 1270 2 83 1301 1 AN2B1S $T=294500 346200 0 0 $X=294500 $Y=345820
X2659 1299 2 1306 1313 1 AN2B1S $T=297600 326040 0 0 $X=297600 $Y=325660
X2660 1279 2 1306 1329 1 AN2B1S $T=301320 326040 0 0 $X=301320 $Y=325660
X2661 1296 2 92 1338 1 AN2B1S $T=303180 305880 0 0 $X=303180 $Y=305500
X2662 1319 2 92 1339 1 AN2B1S $T=303800 315960 1 0 $X=303800 $Y=310540
X2663 1326 2 92 1341 1 AN2B1S $T=305040 265560 1 0 $X=305040 $Y=260140
X2664 1318 2 92 1336 1 AN2B1S $T=305040 275640 1 0 $X=305040 $Y=270220
X2665 1330 2 92 1342 1 AN2B1S $T=305040 285720 0 0 $X=305040 $Y=285340
X2666 260 2 1894 257 1 AN2B1S $T=478640 366360 0 180 $X=475540 $Y=360940
X2667 1901 2 1926 1938 1 AN2B1S $T=487940 326040 0 0 $X=487940 $Y=325660
X2668 1901 2 1964 1960 1 AN2B1S $T=503440 315960 1 180 $X=500340 $Y=315580
X2669 1987 2 2046 2027 1 AN2B1S $T=525140 295800 1 180 $X=522040 $Y=295420
X2670 1987 2 2202 2053 1 AN2B1S $T=562340 285720 0 180 $X=559240 $Y=280300
X2671 2239 2 2425 2437 1 AN2B1S $T=632400 315960 1 180 $X=629300 $Y=315580
X2672 2445 2 2452 2430 1 AN2B1S $T=633640 326040 1 180 $X=630540 $Y=325660
X2673 2445 2 2295 2463 1 AN2B1S $T=633020 346200 1 0 $X=633020 $Y=340780
X2674 2600 2 2609 2622 1 AN2B1S $T=695640 275640 0 0 $X=695640 $Y=275260
X2675 2960 2 2913 2976 1 AN2B1S $T=820260 346200 1 0 $X=820260 $Y=340780
X2676 3329 2 3328 3324 1 AN2B1S $T=979600 285720 0 180 $X=976500 $Y=280300
X2677 3752 2 3754 3758 1 AN2B1S $T=1106080 285720 1 0 $X=1106080 $Y=280300
X2678 1512 1527 1 105 2 1537 OAI12HS $T=365180 295800 1 0 $X=365180 $Y=290380
X2679 178 168 1 10 2 174 OAI12HS $T=401760 265560 0 180 $X=398040 $Y=260140
X2680 263 1914 1 267 2 1925 OAI12HS $T=484220 366360 1 0 $X=484220 $Y=360940
X2681 1956 1951 1 1953 2 1970 OAI12HS $T=499720 346200 1 0 $X=499720 $Y=340780
X2682 1969 1978 1 1962 2 1988 OAI12HS $T=505300 336120 0 0 $X=505300 $Y=335740
X2683 1962 1974 1 1995 2 1985 OAI12HS $T=510880 336120 1 0 $X=510880 $Y=330700
X2684 1981 2056 1 2063 2 2070 OAI12HS $T=525760 326040 0 0 $X=525760 $Y=325660
X2685 2131 2141 1 2143 2 2134 OAI12HS $T=543120 326040 1 0 $X=543120 $Y=320620
X2686 2170 2141 1 2178 2 2172 OAI12HS $T=551180 315960 1 0 $X=551180 $Y=310540
X2687 379 2279 1 386 2 2274 OAI12HS $T=582180 295800 0 0 $X=582180 $Y=295420
X2688 386 2301 1 2310 2 2282 OAI12HS $T=589000 285720 1 0 $X=589000 $Y=280300
X2689 2314 2265 1 2300 2 2289 OAI12HS $T=592720 326040 1 180 $X=589000 $Y=325660
X2690 2288 2309 1 2315 2 2278 OAI12HS $T=590240 336120 0 0 $X=590240 $Y=335740
X2691 2312 2265 1 2319 2 2299 OAI12HS $T=591480 336120 1 0 $X=591480 $Y=330700
X2692 2311 2265 1 2321 2 2298 OAI12HS $T=592100 326040 1 0 $X=592100 $Y=320620
X2693 2334 2309 1 2324 2 2318 OAI12HS $T=598300 336120 1 180 $X=594580 $Y=335740
X2694 2344 2309 1 2328 2 2326 OAI12HS $T=599540 346200 1 180 $X=595820 $Y=345820
X2695 2345 2309 1 2353 2 2356 OAI12HS $T=599540 356280 1 0 $X=599540 $Y=350860
X2696 2330 2363 1 2374 2 2377 OAI12HS $T=606980 326040 0 0 $X=606980 $Y=325660
X2697 2365 2372 1 2378 2 2367 OAI12HS $T=607600 356280 0 0 $X=607600 $Y=355900
X2698 2373 2376 1 2383 2 2362 OAI12HS $T=614420 346200 1 0 $X=614420 $Y=340780
X2699 2378 2398 1 2407 2 2405 OAI12HS $T=616280 356280 0 0 $X=616280 $Y=355900
X2700 2603 2605 1 2587 2 2584 OAI12HS $T=688200 275640 0 0 $X=688200 $Y=275260
X2701 2626 2613 1 2632 2 2636 OAI12HS $T=699360 295800 1 0 $X=699360 $Y=290380
X2702 2638 2652 1 2642 2 2649 OAI12HS $T=708040 315960 0 180 $X=704320 $Y=310540
X2703 2705 2653 1 2720 2 2724 OAI12HS $T=730980 326040 0 180 $X=727260 $Y=320620
X2704 2902 2898 1 2907 2 2913 OAI12HS $T=791740 346200 1 0 $X=791740 $Y=340780
X2705 3524 3506 1 961 2 3488 OAI12HS $T=1040980 265560 0 0 $X=1040980 $Y=265180
X2706 3571 3595 1 3577 2 3599 OAI12HS $T=1062680 315960 0 0 $X=1062680 $Y=315580
X2707 3747 3750 1 3753 2 3614 OAI12HS $T=1104840 305880 0 0 $X=1104840 $Y=305500
X2708 2262 2265 1 2 INV3 $T=582180 336120 0 180 $X=579700 $Y=330700
X2709 2354 2400 1 2 INV3 $T=612560 305880 1 0 $X=612560 $Y=300460
X2710 2381 415 2354 1 2 AN2T $T=610700 326040 0 0 $X=610700 $Y=325660
X2711 2193 1 2203 347 2 ND2P $T=558620 356280 0 0 $X=558620 $Y=355900
X2712 2204 1 2207 349 2 ND2P $T=559860 366360 1 0 $X=559860 $Y=360940
X2713 2240 1 2260 2254 2 ND2P $T=574740 295800 0 0 $X=574740 $Y=295420
X2714 2317 1 2347 2288 2 ND2P $T=598300 336120 1 0 $X=598300 $Y=330700
X2715 2384 1 2355 2283 2 ND2P $T=610700 346200 0 0 $X=610700 $Y=345820
X2716 1112 1102 1119 1 2 1135 HA1 $T=228160 346200 0 0 $X=228160 $Y=345820
X2717 1210 1179 1226 1 2 1233 HA1 $T=261640 326040 0 0 $X=261640 $Y=325660
X2718 1208 1153 1244 1 2 1246 HA1 $T=268460 275640 1 0 $X=268460 $Y=270220
X2719 1165 1238 1276 1 2 1283 HA1 $T=282100 295800 0 0 $X=282100 $Y=295420
X2720 1712 1727 1714 1 2 1711 HA1 $T=421600 295800 1 180 $X=413540 $Y=295420
X2721 1740 1730 207 1 2 1750 HA1 $T=420360 265560 0 0 $X=420360 $Y=265180
X2722 1752 1738 1759 1 2 1775 HA1 $T=425940 346200 1 0 $X=425940 $Y=340780
X2723 1765 1739 1757 1 2 1758 HA1 $T=439580 336120 0 180 $X=431520 $Y=330700
X2724 380 2238 2276 1 2 2287 HA1 $T=576600 275640 1 0 $X=576600 $Y=270220
X2725 2430 2440 2422 1 2 2414 HA1 $T=629300 326040 0 180 $X=621240 $Y=320620
X2726 2463 2491 2506 1 2 2534 HA1 $T=644180 336120 1 0 $X=644180 $Y=330700
X2727 1072 1075 1089 2 1 XOR2HS $T=220720 336120 1 0 $X=220720 $Y=330700
X2728 7 1075 1090 2 1 XOR2HS $T=220720 356280 0 0 $X=220720 $Y=355900
X2729 1094 1073 1103 2 1 XOR2HS $T=225680 285720 1 0 $X=225680 $Y=280300
X2730 1114 1073 1122 2 1 XOR2HS $T=232500 285720 1 0 $X=232500 $Y=280300
X2731 1094 1107 1126 2 1 XOR2HS $T=234360 295800 1 0 $X=234360 $Y=290380
X2732 1117 1107 1130 2 1 XOR2HS $T=234980 305880 0 0 $X=234980 $Y=305500
X2733 1387 97 1400 2 1 XOR2HS $T=318680 356280 1 0 $X=318680 $Y=350860
X2734 1397 1360 1410 2 1 XOR2HS $T=321160 336120 0 0 $X=321160 $Y=335740
X2735 1425 1430 1445 2 1 XOR2HS $T=327360 305880 0 0 $X=327360 $Y=305500
X2736 1442 1452 1458 2 1 XOR2HS $T=331700 265560 0 0 $X=331700 $Y=265180
X2737 1426 1447 1479 2 1 XOR2HS $T=337900 285720 0 0 $X=337900 $Y=285340
X2738 1967 1951 1976 2 1 XOR2HS $T=500960 356280 1 0 $X=500960 $Y=350860
X2739 1980 1978 1990 2 1 XOR2HS $T=505300 346200 0 0 $X=505300 $Y=345820
X2740 2045 2044 2047 2 1 XOR2HS $T=522660 336120 1 0 $X=522660 $Y=330700
X2741 2128 2124 2090 2 1 XOR2HS $T=542500 326040 0 0 $X=542500 $Y=325660
X2742 2156 2141 2111 2 1 XOR2HS $T=548700 326040 0 0 $X=548700 $Y=325660
X2743 2199 2194 2177 2 1 XOR2HS $T=561100 295800 1 180 $X=555520 $Y=295420
X2744 2259 2255 2190 2 1 XOR2HS $T=577220 305880 0 180 $X=571640 $Y=300460
X2745 2267 2265 2242 2 1 XOR2HS $T=579700 326040 1 180 $X=574120 $Y=325660
X2746 2294 2277 2201 2 1 XOR2HS $T=589620 305880 0 180 $X=584040 $Y=300460
X2747 488 482 2621 2 1 XOR2HS $T=695640 265560 0 0 $X=695640 $Y=265180
X2748 2818 2823 2809 2 1 XOR2HS $T=765700 346200 1 180 $X=760120 $Y=345820
X2749 3165 3152 3147 2 1 XOR2HS $T=910160 315960 1 180 $X=904580 $Y=315580
X2750 3239 3237 3200 2 1 XOR2HS $T=938060 305880 0 180 $X=932480 $Y=300460
X2751 3222 3238 3165 2 1 XOR2HS $T=938060 336120 0 180 $X=932480 $Y=330700
X2752 3243 792 3208 2 1 XOR2HS $T=938680 275640 0 0 $X=938680 $Y=275260
X2753 3248 3237 3204 2 1 XOR2HS $T=944880 305880 1 180 $X=939300 $Y=305500
X2754 3249 3237 3159 2 1 XOR2HS $T=944880 336120 0 180 $X=939300 $Y=330700
X2755 3250 3237 3205 2 1 XOR2HS $T=945500 326040 0 180 $X=939920 $Y=320620
X2756 3262 3237 3210 2 1 XOR2HS $T=951700 326040 1 180 $X=946120 $Y=325660
X2757 3263 3237 3238 2 1 XOR2HS $T=951700 336120 0 180 $X=946120 $Y=330700
X2758 2926 2964 2 2951 1 648 MUX2S $T=820880 305880 1 0 $X=820880 $Y=300460
X2759 3018 2964 2 2997 1 660 MUX2S $T=843200 305880 0 180 $X=838860 $Y=300460
X2760 3043 3046 2 3042 1 705 MUX2S $T=858080 295800 0 0 $X=858080 $Y=295420
X2761 497 495 2663 1 2 2689 MAO222 $T=712380 356280 0 0 $X=712380 $Y=355900
X2762 2730 2689 2731 1 2 2734 MAO222 $T=729120 315960 0 0 $X=729120 $Y=315580
X2763 2753 2734 2761 1 2 2782 MAO222 $T=744620 315960 0 0 $X=744620 $Y=315580
X2764 2789 2782 2772 1 2 2802 MAO222 $T=750200 315960 0 0 $X=750200 $Y=315580
X2765 2807 2802 2820 1 2 2831 MAO222 $T=760740 315960 0 0 $X=760740 $Y=315580
X2766 2839 2831 2864 1 2 2847 MAO222 $T=778100 315960 0 180 $X=773140 $Y=310540
X2767 2849 2847 2872 1 2 2859 MAO222 $T=781200 326040 0 180 $X=776240 $Y=320620
X2768 2862 2859 2884 1 2 2877 MAO222 $T=787400 336120 1 180 $X=782440 $Y=335740
X2769 1846 1874 2 1853 1831 1 1900 FA1 $T=461280 285720 1 0 $X=461280 $Y=280300
X2770 1946 1910 2 264 1935 1 1897 FA1 $T=492900 265560 1 180 $X=477400 $Y=265180
X2771 1998 1907 2 1846 1986 1 1947 FA1 $T=511500 295800 0 180 $X=496000 $Y=290380
X2772 1977 1940 2 2021 1984 1 2020 FA1 $T=504680 326040 1 0 $X=504680 $Y=320620
X2773 2038 2054 2 1998 2001 1 2076 FA1 $T=520180 305880 0 0 $X=520180 $Y=305500
X2774 2054 2093 2 2102 1971 1 2086 FA1 $T=525140 295800 0 0 $X=525140 $Y=295420
X2775 2057 2101 2 2108 1982 1 2130 FA1 $T=527000 275640 0 0 $X=527000 $Y=275260
X2776 2068 2037 2 2057 2077 1 2112 FA1 $T=529480 295800 1 0 $X=529480 $Y=290380
X2777 2071 2110 2 321 2083 1 2140 FA1 $T=530100 265560 0 0 $X=530100 $Y=265180
X2778 2083 2130 2 1897 2175 1 338 FA1 $T=536300 265560 1 0 $X=536300 $Y=260140
X2779 2175 353 2 2237 344 1 370 FA1 $T=555520 265560 1 0 $X=555520 $Y=260140
X2780 2333 2375 2 2380 2403 1 2368 FA1 $T=599540 305880 0 0 $X=599540 $Y=305500
X2781 2348 412 2 2386 2357 1 2342 FA1 $T=600160 295800 1 0 $X=600160 $Y=290380
X2782 2320 414 2 2391 416 1 2341 FA1 $T=602020 275640 0 0 $X=602020 $Y=275260
X2783 2357 2387 2 2389 2399 1 2375 FA1 $T=602640 285720 0 0 $X=602640 $Y=285340
X2784 2364 2409 2 2418 2433 1 2395 FA1 $T=608840 315960 1 0 $X=608840 $Y=310540
X2785 433 424 2 2437 2456 1 2416 FA1 $T=636740 265560 0 180 $X=621240 $Y=260140
X2786 2433 2564 2 2471 2557 1 2577 FA1 $T=660920 315960 1 0 $X=660920 $Y=310540
X2787 2599 2525 2 2570 2583 1 2561 FA1 $T=684480 356280 0 180 $X=668980 $Y=350860
X2788 2394 2591 2 2596 2588 1 2415 FA1 $T=673940 336120 1 0 $X=673940 $Y=330700
X2789 2573 2594 2 2338 2606 1 2610 FA1 $T=677660 295800 0 0 $X=677660 $Y=295420
X2790 2401 2586 2 2608 2577 1 2402 FA1 $T=679520 315960 1 0 $X=679520 $Y=310540
X2791 2586 2552 2 2610 2571 1 2591 FA1 $T=682000 305880 0 0 $X=682000 $Y=305500
X2792 2588 2545 2 2599 2598 1 2628 FA1 $T=683860 346200 1 0 $X=683860 $Y=340780
X2793 2441 486 2 2601 2597 1 2447 FA1 $T=685100 356280 0 0 $X=685100 $Y=355900
X2794 2635 484 2 2575 492 1 2601 FA1 $T=702460 366360 0 180 $X=686960 $Y=360940
X2795 2410 2611 2 2612 2628 1 2434 FA1 $T=703080 346200 1 180 $X=687580 $Y=345820
X2796 2611 2561 2 2574 2635 1 2597 FA1 $T=703700 356280 0 180 $X=688200 $Y=350860
X2797 2891 2901 2 2906 2927 1 2895 FA1 $T=802280 295800 0 180 $X=786780 $Y=290380
X2798 2952 2945 2 2946 2958 1 2927 FA1 $T=818400 285720 1 180 $X=802900 $Y=285340
X2799 3035 3019 2 675 3032 1 2958 FA1 $T=854360 285720 0 180 $X=838860 $Y=280300
X2800 378 2 1 382 BUF3 $T=580320 295800 1 0 $X=580320 $Y=290380
X2801 470 2 1 378 BUF3 $T=683240 285720 0 0 $X=683240 $Y=285340
X2802 3089 3068 3081 3083 2 3063 1 AOI13HS $T=874820 326040 0 180 $X=871100 $Y=320620
X2803 3619 3631 3629 3624 2 3621 1 AOI13HS $T=1073840 295800 0 180 $X=1070120 $Y=290380
X2804 3779 3772 3776 3743 2 3705 1 AOI13HS $T=1114760 295800 0 180 $X=1111040 $Y=290380
X2805 1464 1 2 1472 1484 1461 1070 ICV_27 $T=336660 315960 1 0 $X=336660 $Y=310540
X2806 112 1 2 120 1504 1509 1070 ICV_27 $T=345340 265560 0 0 $X=345340 $Y=265180
X2807 2669 1 2 2664 2647 2696 1070 ICV_27 $T=709280 295800 1 0 $X=709280 $Y=290380
X2808 642 1 2 650 652 656 1070 ICV_27 $T=824600 326040 0 0 $X=824600 $Y=325660
X2809 3147 1 2 3146 3154 3166 1070 ICV_27 $T=900240 265560 0 0 $X=900240 $Y=265180
X2810 750 1 2 3183 757 762 1070 ICV_27 $T=910780 295800 1 0 $X=910780 $Y=290380
X2811 3186 1 2 3175 3199 3181 1070 ICV_27 $T=917600 265560 1 0 $X=917600 $Y=260140
X2812 768 1 2 3219 778 783 1070 ICV_27 $T=925040 295800 1 0 $X=925040 $Y=290380
X2813 774 1 2 3223 3229 3232 1070 ICV_27 $T=928140 265560 1 0 $X=928140 $Y=260140
X2814 787 1 2 3246 800 809 1070 ICV_27 $T=941160 285720 0 0 $X=941160 $Y=285340
X2815 804 1 2 816 803 3265 1070 ICV_27 $T=949840 265560 1 0 $X=949840 $Y=260140
X2816 818 1 2 824 825 834 1070 ICV_27 $T=954180 295800 1 0 $X=954180 $Y=290380
X2817 3272 1 2 3275 829 835 1070 ICV_27 $T=956660 315960 1 0 $X=956660 $Y=310540
X2818 837 1 2 843 844 850 1070 ICV_27 $T=966580 315960 1 0 $X=966580 $Y=310540
X2819 842 1 2 848 849 855 1070 ICV_27 $T=970300 305880 0 0 $X=970300 $Y=305500
X2820 858 1 2 866 868 875 1070 ICV_27 $T=981460 305880 0 0 $X=981460 $Y=305500
X2821 883 1 2 890 3365 3377 1070 ICV_27 $T=993860 326040 1 0 $X=993860 $Y=320620
X2822 908 1 2 912 914 919 1070 ICV_27 $T=1011840 336120 1 0 $X=1011840 $Y=330700
X2823 3441 1 2 3455 921 935 1070 ICV_27 $T=1019900 315960 0 0 $X=1019900 $Y=315580
X2824 920 1 2 923 926 936 1070 ICV_27 $T=1021140 336120 0 0 $X=1021140 $Y=335740
X2825 940 1 2 946 947 3467 1070 ICV_27 $T=1031060 336120 0 0 $X=1031060 $Y=335740
X2826 967 1 2 976 952 3552 1070 ICV_27 $T=1044700 346200 0 0 $X=1044700 $Y=345820
X2827 969 1 2 977 978 987 1070 ICV_27 $T=1045320 336120 0 0 $X=1045320 $Y=335740
X2828 1044 1 2 1047 1048 1052 1070 ICV_27 $T=1116000 346200 1 0 $X=1116000 $Y=340780
X2829 1912 1887 1 2 BUF6 $T=491660 295800 0 0 $X=491660 $Y=295420
X2830 281 1912 1 2 BUF6 $T=498480 265560 1 0 $X=498480 $Y=260140
X2831 1420 104 1334 1437 2 1 MXL2HS $T=334800 356280 0 180 $X=329220 $Y=350860
X2832 1436 104 1324 1463 2 1 MXL2HS $T=331700 346200 0 0 $X=331700 $Y=345820
X2833 1409 104 1368 1475 2 1 MXL2HS $T=334800 336120 0 0 $X=334800 $Y=335740
X2834 1462 1457 1381 1474 2 1 MXL2HS $T=342860 315960 1 180 $X=337280 $Y=315580
X2835 1448 1457 1383 1491 2 1 MXL2HS $T=339760 285720 1 0 $X=339760 $Y=280300
X2836 1487 1457 1449 1497 2 1 MXL2HS $T=341620 275640 0 0 $X=341620 $Y=275260
X2837 1464 1457 1444 1503 2 1 MXL2HS $T=344720 285720 0 0 $X=344720 $Y=285340
X2838 1484 1457 1441 1511 2 1 MXL2HS $T=345960 315960 0 0 $X=345960 $Y=315580
X2839 1504 130 1398 1531 2 1 MXL2HS $T=353400 265560 1 0 $X=353400 $Y=260140
X2840 1075 12 1100 1099 1 2 HA1P $T=220720 356280 1 0 $X=220720 $Y=350860
X2841 1107 1106 1088 1084 1 2 HA1P $T=231880 295800 1 180 $X=222580 $Y=295420
X2842 1094 1088 1097 1086 1 2 HA1P $T=234360 285720 1 180 $X=225060 $Y=285340
X2843 1073 1097 22 1093 1 2 HA1P $T=226300 265560 0 0 $X=226300 $Y=265180
X2844 1117 1100 1106 1098 1 2 HA1P $T=237460 315960 1 180 $X=228160 $Y=315580
X2845 2745 532 2756 2760 1 2 HA1P $T=736560 356280 0 0 $X=736560 $Y=355900
X2846 2749 2756 2758 2766 1 2 HA1P $T=737180 346200 0 0 $X=737180 $Y=345820
X2847 2728 2758 2770 2777 1 2 HA1P $T=738420 336120 0 0 $X=738420 $Y=335740
X2848 2786 2770 2803 2812 1 2 HA1P $T=748340 346200 1 0 $X=748340 $Y=340780
X2849 2791 2803 2837 2825 1 2 HA1P $T=759500 346200 1 0 $X=759500 $Y=340780
X2850 2841 2837 2863 2846 1 2 HA1P $T=770660 346200 1 0 $X=770660 $Y=340780
X2851 2840 2863 2823 2843 1 2 HA1P $T=783060 346200 1 180 $X=773760 $Y=345820
X2852 2270 385 1 2275 2 AN2S $T=585280 336120 0 180 $X=582800 $Y=330700
X2853 2166 2179 1 2164 339 2160 2 OAI22H $T=556760 265560 1 180 $X=549320 $Y=265180
X2854 2326 365 2304 1 2 XNR2H $T=598300 356280 1 180 $X=589620 $Y=355900
X2855 1361 1367 2 1360 1350 1 AOI12H $T=316820 336120 1 180 $X=310620 $Y=335740
X2856 1423 1427 2 1430 1419 1 AOI12H $T=326120 315960 0 0 $X=326120 $Y=315580
X2857 1408 1451 2 1447 1422 1 AOI12H $T=334800 295800 0 180 $X=328600 $Y=290380
X2858 1434 1453 2 1452 1440 1 AOI12H $T=331700 275640 1 0 $X=331700 $Y=270220
X2859 2148 2144 2 2178 2153 1 AOI12H $T=547460 305880 0 0 $X=547460 $Y=305500
X2860 2384 2362 2 2297 2405 1 AOI12H $T=613800 356280 1 0 $X=613800 $Y=350860
X2861 3733 3732 2 3666 1 3727 AN3B2S $T=1103600 315960 0 180 $X=1099880 $Y=310540
X2862 3775 3627 2 3753 1 3783 AN3B2S $T=1112280 326040 1 0 $X=1112280 $Y=320620
X2863 892 3354 3425 2 1 904 OR3 $T=1006260 265560 1 0 $X=1006260 $Y=260140
X2864 1902 1888 1 2 INV2CK $T=479260 275640 0 180 $X=476780 $Y=270220
X2865 3046 2982 1 2 INV2CK $T=863040 295800 0 0 $X=863040 $Y=295420
X2866 2623 2719 1 2694 505 2663 2 MOAI1HT $T=730360 285720 1 180 $X=711760 $Y=285340
X2867 2623 2779 1 2694 531 2731 2 MOAI1HT $T=750820 295800 0 180 $X=732220 $Y=290380
X2868 2942 2924 1 2917 603 2884 2 MOAI1HT $T=807240 336120 1 180 $X=788640 $Y=335740
X2869 2623 2926 1 2917 2954 2872 2 MOAI1HT $T=816540 305880 0 180 $X=797940 $Y=300460
X2870 2942 2962 1 2917 627 2948 2 MOAI1HT $T=824600 326040 1 180 $X=806000 $Y=325660
X2871 2942 2885 1 2917 641 2981 2 MOAI1HT $T=811580 336120 0 0 $X=811580 $Y=335740
X2872 3004 3002 1 2972 654 2761 2 MOAI1HT $T=837620 295800 0 180 $X=819020 $Y=290380
X2873 2942 2844 1 2972 668 3001 2 MOAI1HT $T=828320 336120 1 0 $X=828320 $Y=330700
X2874 3004 2985 1 2972 678 3031 2 MOAI1HT $T=833280 336120 0 0 $X=833280 $Y=335740
X2875 3004 3038 1 2972 682 2772 2 MOAI1HT $T=858700 285720 1 180 $X=840100 $Y=285340
X2876 3004 3043 1 2972 689 2820 2 MOAI1HT $T=858700 295800 0 180 $X=840100 $Y=290380
X2877 3004 3018 1 2972 685 2864 2 MOAI1HT $T=859320 315960 1 180 $X=840720 $Y=315580
X2878 2639 2623 1 2 2694 OR2B1 $T=723540 305880 0 0 $X=723540 $Y=305500
X2879 2639 2617 1 2620 489 2 2613 2630 493 OAI222S $T=704940 295800 1 180 $X=699360 $Y=295420
X2880 2639 2623 1 490 2 OR2T $T=704320 315960 0 180 $X=698120 $Y=310540
X2881 2157 2184 2 2215 2191 1 AOI12HP $T=553660 305880 0 0 $X=553660 $Y=305500
X2882 2262 2271 2 383 2284 1 AOI12HP $T=575980 356280 1 0 $X=575980 $Y=350860
X2883 2250 2260 2 2281 2282 1 AOI12HP $T=576600 285720 0 0 $X=576600 $Y=285340
X2884 2271 2262 2 390 2284 1 AOI12HP $T=579080 346200 0 0 $X=579080 $Y=345820
X2885 2337 2347 2 2315 2377 1 AOI12HP $T=602020 336120 1 0 $X=602020 $Y=330700
X2886 1401 1360 1 1384 1427 2 OAI12H $T=323020 326040 0 0 $X=323020 $Y=325660
X2887 1405 1430 1 1403 1451 2 OAI12H $T=326740 305880 1 0 $X=326740 $Y=300460
X2888 1429 1452 1 1443 106 2 OAI12H $T=331080 265560 1 0 $X=331080 $Y=260140
X2889 2118 2097 1 2116 2157 2 OAI12H $T=543120 315960 0 0 $X=543120 $Y=315580
X2890 333 2178 1 340 2191 2 OAI12H $T=552420 305880 1 0 $X=552420 $Y=300460
X2891 2233 357 1 352 2250 2 OAI12H $T=569780 285720 0 0 $X=569780 $Y=285340
X2892 2321 2329 1 2336 2337 2 OAI12H $T=598920 315960 0 0 $X=598920 $Y=315580
X2893 1352 97 1 1364 1367 2 OAI12HP $T=308140 356280 1 0 $X=308140 $Y=350860
X2894 1421 1447 1 1411 1453 2 OAI12HP $T=327360 285720 0 0 $X=327360 $Y=285340
X2895 2283 2315 1 2297 2284 2 OAI12HP $T=597680 356280 0 180 $X=587140 $Y=350860
X2896 2271 2288 1 2283 2 NR2T $T=582800 346200 1 0 $X=582800 $Y=340780
X2897 2254 2215 1 2281 2262 2 OAI12HT $T=572260 305880 0 0 $X=572260 $Y=305500
.ENDS
***************************************
.SUBCKT TIE1 O VCC GND
** N=4 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT TIE0 O VCC GND
** N=4 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DELC I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA13S B3 B2 B1 A1 GND VCC O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_33 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 186 187 188 189 190 191 192 193 194 196 197 198 199 200 201 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223
+ 224 225 226 228 229 230 231 232 233 234 235 236 237 238 240 241 242 243 244 245
+ 246 247 248 250 251 252 253 254 255 256 257 258 259 260 261 263 264 265 266 267
+ 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283 284 285 286 287
+ 288 289 290 291 292 293 294 295 296 297 298 299 300 301 302 303 304 305 306 307
+ 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324 325 326 327
+ 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347
+ 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362 363 364 365 366 367
+ 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382 383 384 385 386 387
+ 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406 407
+ 408 421 435
** N=1297 EP=403 IP=5770 FDC=0
X0 408 407 407 407 421 407 405 YA2GSD $T=1349740 190760 0 90 $X=1210240 $Y=193610
X1 441 2 439 1 INV1S $T=223200 245400 1 180 $X=221960 $Y=245020
X2 447 2 446 1 INV1S $T=229400 245400 1 180 $X=228160 $Y=245020
X3 452 2 453 1 INV1S $T=233740 235320 1 0 $X=233740 $Y=229900
X4 459 2 460 1 INV1S $T=248000 235320 0 0 $X=248000 $Y=234940
X5 18 2 464 1 INV1S $T=249240 235320 0 0 $X=249240 $Y=234940
X6 16 2 22 1 INV1S $T=249860 255480 0 0 $X=249860 $Y=255100
X7 24 2 469 1 INV1S $T=256680 235320 0 0 $X=256680 $Y=234940
X8 463 2 28 1 INV1S $T=258540 235320 1 0 $X=258540 $Y=229900
X9 26 2 473 1 INV1S $T=258540 235320 0 0 $X=258540 $Y=234940
X10 17 2 475 1 INV1S $T=260400 235320 1 0 $X=260400 $Y=229900
X11 460 2 34 1 INV1S $T=265360 235320 0 0 $X=265360 $Y=234940
X12 34 2 480 1 INV1S $T=266600 255480 0 180 $X=265360 $Y=250060
X13 27 2 483 1 INV1S $T=266600 255480 1 0 $X=266600 $Y=250060
X14 487 2 493 1 INV1S $T=275900 225240 0 0 $X=275900 $Y=224860
X15 485 2 495 1 INV1S $T=275900 235320 0 0 $X=275900 $Y=234940
X16 488 2 494 1 INV1S $T=277760 245400 0 0 $X=277760 $Y=245020
X17 549 2 550 1 INV1S $T=328600 255480 1 0 $X=328600 $Y=250060
X18 563 2 566 1 INV1S $T=339140 255480 1 0 $X=339140 $Y=250060
X19 567 2 575 1 INV1S $T=345340 235320 1 0 $X=345340 $Y=229900
X20 577 2 578 1 INV1S $T=346580 225240 0 0 $X=346580 $Y=224860
X21 608 2 612 1 INV1S $T=384400 235320 0 180 $X=383160 $Y=229900
X22 74 2 69 1 INV1S $T=391220 245400 1 180 $X=389980 $Y=245020
X23 76 2 72 1 INV1S $T=393700 255480 1 180 $X=392460 $Y=255100
X24 78 2 609 1 INV1S $T=395560 255480 1 180 $X=394320 $Y=255100
X25 81 2 82 1 INV1S $T=400520 255480 0 0 $X=400520 $Y=255100
X26 83 2 74 1 INV1S $T=403000 255480 1 180 $X=401760 $Y=255100
X27 597 2 79 1 INV1S $T=403620 235320 1 180 $X=402380 $Y=234940
X28 625 2 83 1 INV1S $T=404860 255480 1 180 $X=403620 $Y=255100
X29 627 2 626 1 INV1S $T=406100 235320 0 180 $X=404860 $Y=229900
X30 597 2 628 1 INV1S $T=404860 235320 0 0 $X=404860 $Y=234940
X31 626 2 631 1 INV1S $T=406100 235320 1 0 $X=406100 $Y=229900
X32 631 2 637 1 INV1S $T=408580 235320 1 0 $X=408580 $Y=229900
X33 624 2 629 1 INV1S $T=408580 255480 0 0 $X=408580 $Y=255100
X34 101 2 99 1 INV1S $T=446400 245400 0 180 $X=445160 $Y=239980
X35 101 2 100 1 INV1S $T=445160 255480 0 0 $X=445160 $Y=255100
X36 117 2 680 1 INV1S $T=481120 255480 0 180 $X=479880 $Y=250060
X37 117 2 687 1 INV1S $T=481740 255480 1 0 $X=481740 $Y=250060
X38 741 2 753 1 INV1S $T=574120 255480 0 0 $X=574120 $Y=255100
X39 811 2 816 1 INV1S $T=672080 255480 0 180 $X=670840 $Y=250060
X40 825 2 831 1 INV1S $T=691920 245400 1 0 $X=691920 $Y=239980
X41 835 2 843 1 INV1S $T=698740 235320 0 0 $X=698740 $Y=234940
X42 839 2 208 1 INV1S $T=700600 255480 0 180 $X=699360 $Y=250060
X43 826 2 842 1 INV1S $T=700600 245400 1 0 $X=700600 $Y=239980
X44 211 2 210 1 INV1S $T=702460 255480 0 0 $X=702460 $Y=255100
X45 850 2 845 1 INV1S $T=706800 245400 0 180 $X=705560 $Y=239980
X46 212 2 850 1 INV1S $T=705560 255480 0 0 $X=705560 $Y=255100
X47 850 2 853 1 INV1S $T=708040 235320 0 0 $X=708040 $Y=234940
X48 858 2 861 1 INV1S $T=713000 235320 0 0 $X=713000 $Y=234940
X49 869 2 868 1 INV1S $T=717340 235320 0 0 $X=717340 $Y=234940
X50 870 2 859 1 INV1S $T=719820 255480 0 180 $X=718580 $Y=250060
X51 252 2 940 1 INV1S $T=787400 255480 1 180 $X=786160 $Y=255100
X52 256 2 888 1 INV1S $T=791120 255480 1 0 $X=791120 $Y=250060
X53 258 2 942 1 INV1S $T=796080 255480 1 180 $X=794840 $Y=255100
X54 265 2 909 1 INV1S $T=797940 255480 0 180 $X=796700 $Y=250060
X55 268 2 966 1 INV1S $T=818400 255480 0 180 $X=817160 $Y=250060
X56 270 2 896 1 INV1S $T=819640 245400 1 180 $X=818400 $Y=245020
X57 276 2 977 1 INV1S $T=827080 255480 0 0 $X=827080 $Y=255100
X58 283 2 996 1 INV1S $T=839480 255480 1 0 $X=839480 $Y=250060
X59 286 2 985 1 INV1S $T=845060 245400 1 180 $X=843820 $Y=245020
X60 292 2 992 1 INV1S $T=859940 245400 1 0 $X=859940 $Y=239980
X61 1022 2 278 1 INV1S $T=866140 245400 1 180 $X=864900 $Y=245020
X62 287 2 296 1 INV1S $T=872960 255480 0 0 $X=872960 $Y=255100
X63 297 2 987 1 INV1S $T=876060 235320 0 180 $X=874820 $Y=229900
X64 1034 2 998 1 INV1S $T=879160 245400 1 180 $X=877920 $Y=245020
X65 1037 2 1004 1 INV1S $T=882260 235320 0 180 $X=881020 $Y=229900
X66 299 2 1039 1 INV1S $T=884740 245400 1 180 $X=883500 $Y=245020
X67 1048 2 1013 1 INV1S $T=886600 235320 1 180 $X=885360 $Y=234940
X68 1052 2 1007 1 INV1S $T=890320 245400 0 180 $X=889080 $Y=239980
X69 1063 2 1058 1 INV1S $T=897760 255480 0 180 $X=896520 $Y=250060
X70 1098 2 1090 1 INV1S $T=941780 245400 1 180 $X=940540 $Y=245020
X71 310 2 1098 1 INV1S $T=947980 245400 0 0 $X=947980 $Y=245020
X72 1098 2 1105 1 INV1S $T=949840 245400 1 0 $X=949840 $Y=239980
X73 327 2 338 1 INV1S $T=991380 255480 1 0 $X=991380 $Y=250060
X74 323 2 341 1 INV1S $T=996340 255480 0 0 $X=996340 $Y=255100
X75 1147 2 1152 1 INV1S $T=1017420 225240 1 180 $X=1016180 $Y=224860
X76 1155 2 1169 1 INV1S $T=1024240 235320 0 0 $X=1024240 $Y=234940
X77 1179 2 1188 1 INV1S $T=1037260 225240 1 180 $X=1036020 $Y=224860
X78 1191 2 1179 1 INV1S $T=1038500 225240 1 180 $X=1037260 $Y=224860
X79 366 2 1191 1 INV1S $T=1039120 235320 1 180 $X=1037880 $Y=234940
X80 363 2 1167 1 INV1S $T=1038500 245400 0 0 $X=1038500 $Y=245020
X81 1194 2 355 1 INV1S $T=1039740 255480 0 180 $X=1038500 $Y=250060
X82 1191 2 1196 1 INV1S $T=1039740 225240 0 0 $X=1039740 $Y=224860
X83 1186 2 364 1 INV1S $T=1042840 255480 0 180 $X=1041600 $Y=250060
X84 372 2 370 1 INV1S $T=1045320 255480 0 180 $X=1044080 $Y=250060
X85 1178 2 1204 1 INV1S $T=1049660 225240 1 180 $X=1048420 $Y=224860
X86 1213 2 1168 1 INV1S $T=1050900 235320 1 180 $X=1049660 $Y=234940
X87 1213 2 1212 1 INV1S $T=1050900 245400 1 180 $X=1049660 $Y=245020
X88 373 2 1216 1 INV1S $T=1051520 245400 0 0 $X=1051520 $Y=245020
X89 353 2 362 1 INV1S $T=1054620 255480 0 0 $X=1054620 $Y=255100
X90 1219 2 1223 1 INV1S $T=1057100 245400 0 0 $X=1057100 $Y=245020
X91 1223 2 1160 1 INV1S $T=1060200 245400 1 180 $X=1058960 $Y=245020
X92 365 2 1222 1 INV1S $T=1064540 245400 0 180 $X=1063300 $Y=239980
X93 1225 2 1176 1 INV1S $T=1065780 245400 1 0 $X=1065780 $Y=239980
X94 1223 2 1234 1 INV1S $T=1067020 235320 0 0 $X=1067020 $Y=234940
X95 377 2 1238 1 INV1S $T=1068260 245400 1 0 $X=1068260 $Y=239980
X96 387 2 1213 1 INV1S $T=1071980 255480 0 180 $X=1070740 $Y=250060
X97 1241 2 385 1 INV1S $T=1073220 245400 0 0 $X=1073220 $Y=245020
X98 384 2 387 1 INV1S $T=1073840 255480 0 0 $X=1073840 $Y=255100
X99 388 2 1189 1 INV1S $T=1077560 245400 1 0 $X=1077560 $Y=239980
X100 1235 2 1161 1 INV1S $T=1077560 245400 0 0 $X=1077560 $Y=245020
X101 1259 2 1260 1 INV1S $T=1094920 235320 1 0 $X=1094920 $Y=229900
X102 1274 2 1271 1 INV1S $T=1102980 235320 0 0 $X=1102980 $Y=234940
X103 1282 2 1284 1 INV1S $T=1106700 255480 1 0 $X=1106700 $Y=250060
X104 1280 2 1285 1 INV1S $T=1109180 235320 0 0 $X=1109180 $Y=234940
X105 1278 2 1288 1 INV1S $T=1111660 245400 0 0 $X=1111660 $Y=245020
X106 1295 2 1289 1 INV1S $T=1121580 255480 1 180 $X=1120340 $Y=255100
X107 3 1 2 4 BUF1S $T=223200 225240 0 180 $X=220720 $Y=219820
X108 450 1 2 441 BUF1S $T=233120 255480 1 0 $X=233120 $Y=250060
X109 452 1 2 463 BUF1S $T=245520 235320 1 0 $X=245520 $Y=229900
X110 463 1 2 25 BUF1S $T=251720 245400 1 0 $X=251720 $Y=239980
X111 461 1 2 31 BUF1S $T=260400 245400 0 0 $X=260400 $Y=245020
X112 20 1 2 481 BUF1S $T=266600 245400 0 0 $X=266600 $Y=245020
X113 33 1 2 484 BUF1S $T=274040 255480 1 0 $X=274040 $Y=250060
X114 46 1 2 512 BUF1S $T=307520 255480 0 0 $X=307520 $Y=255100
X115 52 1 2 3 BUF1S $T=329840 225240 0 180 $X=327360 $Y=219820
X116 62 1 2 594 BUF1S $T=357740 235320 0 0 $X=357740 $Y=234940
X117 63 1 2 602 BUF1S $T=369520 245400 0 0 $X=369520 $Y=245020
X118 73 1 2 608 BUF1S $T=391840 225240 1 180 $X=389360 $Y=224860
X119 72 1 2 617 BUF1S $T=389360 255480 1 0 $X=389360 $Y=250060
X120 619 1 2 68 BUF1S $T=397420 235320 0 180 $X=394940 $Y=229900
X121 79 1 2 619 BUF1S $T=400520 235320 0 180 $X=398040 $Y=229900
X122 639 1 2 643 BUF1S $T=414160 235320 1 0 $X=414160 $Y=229900
X123 151 1 2 761 BUF1S $T=582800 255480 0 0 $X=582800 $Y=255100
X124 822 1 2 823 BUF1S $T=677660 235320 1 0 $X=677660 $Y=229900
X125 217 1 2 851 BUF1S $T=716720 245400 0 180 $X=714240 $Y=239980
X126 888 1 2 963 BUF1S $T=808480 235320 0 0 $X=808480 $Y=234940
X127 966 1 2 893 BUF1S $T=814680 255480 0 180 $X=812200 $Y=250060
X128 274 1 2 890 BUF1S $T=825220 245400 1 180 $X=822740 $Y=245020
X129 977 1 2 894 BUF1S $T=826460 245400 0 180 $X=823980 $Y=239980
X130 278 1 2 898 BUF1S $T=831420 245400 0 180 $X=828940 $Y=239980
X131 985 1 2 902 BUF1S $T=833900 245400 1 180 $X=831420 $Y=245020
X132 987 1 2 936 BUF1S $T=834520 245400 0 180 $X=832040 $Y=239980
X133 992 1 2 912 BUF1S $T=839480 245400 1 180 $X=837000 $Y=245020
X134 996 1 2 907 BUF1S $T=843200 245400 1 180 $X=840720 $Y=245020
X135 998 1 2 905 BUF1S $T=846300 255480 0 180 $X=843820 $Y=250060
X136 287 1 2 945 BUF1S $T=848160 245400 1 180 $X=845680 $Y=245020
X137 1007 1 2 934 BUF1S $T=851880 245400 1 180 $X=849400 $Y=245020
X138 1004 1 2 955 BUF1S $T=851260 235320 0 0 $X=851260 $Y=234940
X139 1013 1 2 929 BUF1S $T=857460 235320 1 180 $X=854980 $Y=234940
X140 312 1 2 315 BUF1S $T=923800 255480 1 0 $X=923800 $Y=250060
X141 1091 1 2 1078 BUF1S $T=938060 255480 0 0 $X=938060 $Y=255100
X142 1101 1 2 319 BUF1S $T=947980 235320 0 180 $X=945500 $Y=229900
X143 345 1 2 302 BUF1S $T=1003160 225240 0 180 $X=1000680 $Y=219820
X144 1167 1 2 1208 BUF1S $T=1044700 245400 0 0 $X=1044700 $Y=245020
X145 375 1 2 1187 BUF1S $T=1050900 255480 1 180 $X=1048420 $Y=255100
X146 374 1 2 1224 BUF1S $T=1060200 245400 0 0 $X=1060200 $Y=245020
X147 386 1 2 1192 BUF1S $T=1077560 235320 0 180 $X=1075080 $Y=229900
X148 1245 1 2 1235 BUF1S $T=1075080 245400 1 0 $X=1075080 $Y=239980
X149 1165 1 2 1241 BUF1S $T=1075080 245400 0 0 $X=1075080 $Y=245020
X150 393 1 2 1251 BUF1S $T=1095540 245400 0 180 $X=1093060 $Y=239980
X151 394 1 2 393 BUF1S $T=1100500 255480 1 180 $X=1098020 $Y=255100
X152 1266 1 2 1267 BUF1S $T=1098640 255480 1 0 $X=1098640 $Y=250060
X153 404 1 2 345 BUF1S $T=1112900 225240 0 180 $X=1110420 $Y=219820
X154 5 1 2 9 DELB $T=222580 255480 1 0 $X=222580 $Y=250060
X155 446 1 2 443 DELB $T=227540 255480 1 0 $X=227540 $Y=250060
X156 451 1 2 452 DELB $T=233740 225240 0 0 $X=233740 $Y=224860
X157 12 1 2 14 DELB $T=236220 255480 1 0 $X=236220 $Y=250060
X158 640 1 2 597 DELB $T=412920 225240 0 0 $X=412920 $Y=224860
X159 642 1 2 625 DELB $T=414780 245400 1 0 $X=414780 $Y=239980
X160 817 1 2 818 DELB $T=671460 245400 1 0 $X=671460 $Y=239980
X161 821 1 2 820 DELB $T=676420 245400 1 0 $X=676420 $Y=239980
X162 857 1 2 865 DELB $T=709900 245400 0 0 $X=709900 $Y=245020
X163 860 1 2 869 DELB $T=713620 235320 1 0 $X=713620 $Y=229900
X164 871 1 2 876 DELB $T=720440 255480 1 0 $X=720440 $Y=250060
X165 877 1 2 879 DELB $T=741520 235320 0 0 $X=741520 $Y=234940
X166 1070 1 2 1071 DELB $T=915740 235320 0 0 $X=915740 $Y=234940
X167 1254 1 2 1259 DELB $T=1086240 235320 1 0 $X=1086240 $Y=229900
X168 1296 1 2 1295 DELB $T=1124680 255480 0 0 $X=1124680 $Y=255100
X169 51 1 2 555 DELA $T=331080 255480 0 0 $X=331080 $Y=255100
X170 61 1 2 600 DELA $T=365800 235320 1 0 $X=365800 $Y=229900
X171 621 1 2 618 DELA $T=396800 245400 1 0 $X=396800 $Y=239980
X172 824 1 2 819 DELA $T=681380 245400 1 0 $X=681380 $Y=239980
X173 843 1 2 844 DELA $T=701220 225240 1 0 $X=701220 $Y=219820
X174 221 1 2 223 DELA $T=725400 255480 1 0 $X=725400 $Y=250060
X175 1065 1 2 1067 DELA $T=907680 245400 0 0 $X=907680 $Y=245020
X176 1068 1 2 1069 DELA $T=913880 235320 1 0 $X=913880 $Y=229900
X177 1074 1 2 1073 DELA $T=920700 225240 1 0 $X=920700 $Y=219820
X178 1075 1 2 1077 DELA $T=923800 235320 0 0 $X=923800 $Y=234940
X179 1088 1 2 1072 DELA $T=931240 235320 0 0 $X=931240 $Y=234940
X180 1095 1 2 1089 DELA $T=939300 235320 0 0 $X=939300 $Y=234940
X181 1096 1 2 1086 DELA $T=941780 245400 1 0 $X=941780 $Y=239980
X182 1246 1 2 1252 DELA $T=1080040 235320 1 0 $X=1080040 $Y=229900
X183 1279 1 2 1287 DELA $T=1106700 245400 0 0 $X=1106700 $Y=245020
X184 1292 1 2 1281 DELA $T=1116620 235320 0 0 $X=1116620 $Y=234940
X185 437 6 10 2 1 447 QDFFRBN $T=220720 255480 0 0 $X=220720 $Y=255100
X186 438 6 10 2 1 450 QDFFRBN $T=221340 235320 0 0 $X=221340 $Y=234940
X187 440 6 10 2 1 451 QDFFRBN $T=221960 225240 0 0 $X=221960 $Y=224860
X188 586 6 63 2 1 58 QDFFRBN $T=367040 255480 1 180 $X=355260 $Y=255100
X189 589 6 63 2 1 62 QDFFRBN $T=368280 255480 0 180 $X=356500 $Y=250060
X190 599 6 602 2 1 61 QDFFRBN $T=380060 245400 0 180 $X=368280 $Y=239980
X191 618 6 602 2 1 76 QDFFRBN $T=392460 245400 0 0 $X=392460 $Y=245020
X192 645 6 602 2 1 642 QDFFRBN $T=426560 245400 1 180 $X=414780 $Y=245020
X193 86 6 602 2 1 85 QDFFRBN $T=427180 255480 1 180 $X=415400 $Y=255100
X194 643 6 602 2 1 627 QDFFRBN $T=430280 235320 0 180 $X=418500 $Y=229900
X195 644 6 602 2 1 640 QDFFRBN $T=430280 235320 1 180 $X=418500 $Y=234940
X196 818 199 201 2 1 825 QDFFRBN $T=675180 245400 0 0 $X=675180 $Y=245020
X197 819 199 201 2 1 826 QDFFRBN $T=675180 255480 1 0 $X=675180 $Y=250060
X198 820 199 201 2 1 827 QDFFRBN $T=675800 235320 0 0 $X=675800 $Y=234940
X199 200 199 201 2 1 205 QDFFRBN $T=679520 255480 0 0 $X=679520 $Y=255100
X200 823 199 201 2 1 835 QDFFRBN $T=680140 235320 1 0 $X=680140 $Y=229900
X201 865 199 220 2 1 870 QDFFRBN $T=730980 245400 1 180 $X=719200 $Y=245020
X202 222 199 220 2 1 219 QDFFRBN $T=731600 255480 1 180 $X=719820 $Y=255100
X203 876 199 220 2 1 854 QDFFRBN $T=734080 245400 0 180 $X=722300 $Y=239980
X204 873 199 220 2 1 860 QDFFRBN $T=737180 235320 0 180 $X=725400 $Y=229900
X205 879 199 220 2 1 874 QDFFRBN $T=741520 235320 1 180 $X=729740 $Y=234940
X206 1071 308 306 2 1 1034 QDFFRBN $T=912640 245400 0 180 $X=900860 $Y=239980
X207 1069 308 306 2 1 1048 QDFFRBN $T=915740 235320 1 180 $X=903960 $Y=234940
X208 1073 308 306 2 1 1052 QDFFRBN $T=916360 225240 0 180 $X=904580 $Y=219820
X209 1067 308 306 2 1 1022 QDFFRBN $T=916360 255480 0 180 $X=904580 $Y=250060
X210 1072 308 306 2 1 1037 QDFFRBN $T=919460 225240 1 180 $X=907680 $Y=224860
X211 1066 308 310 2 1 1075 QDFFRBN $T=911400 255480 0 0 $X=911400 $Y=255100
X212 316 308 1090 2 1 1091 QDFFRBN $T=926280 255480 0 0 $X=926280 $Y=255100
X213 1081 308 1090 2 1 1096 QDFFRBN $T=926900 245400 0 0 $X=926900 $Y=245020
X214 1087 308 1090 2 1 1095 QDFFRBN $T=930000 245400 1 0 $X=930000 $Y=239980
X215 1093 308 310 2 1 323 QDFFRBN $T=938060 255480 1 0 $X=938060 $Y=250060
X216 1108 308 310 2 1 1100 QDFFRBN $T=964720 255480 0 180 $X=952940 $Y=250060
X217 1110 308 1105 2 1 1102 QDFFRBN $T=965340 235320 1 180 $X=953560 $Y=234940
X218 1099 308 1105 2 1 327 QDFFRBN $T=953560 245400 0 0 $X=953560 $Y=245020
X219 1122 308 1105 2 1 1097 QDFFRBN $T=965960 225240 1 180 $X=954180 $Y=224860
X220 1111 308 1105 2 1 1104 QDFFRBN $T=967820 235320 0 180 $X=956040 $Y=229900
X221 1137 308 1105 2 1 1103 QDFFRBN $T=980840 225240 0 180 $X=969060 $Y=219820
X222 1158 308 350 2 1 1101 QDFFRBN $T=1023000 245400 0 180 $X=1011220 $Y=239980
X223 1161 308 350 2 1 1150 QDFFRBN $T=1024860 255480 0 180 $X=1013080 $Y=250060
X224 1255 391 390 2 1 1246 QDFFRBN $T=1091820 225240 1 180 $X=1080040 $Y=224860
X225 1258 391 390 2 1 1245 QDFFRBN $T=1091820 245400 0 180 $X=1080040 $Y=239980
X226 392 391 390 2 1 1248 QDFFRBN $T=1093680 255480 1 180 $X=1081900 $Y=255100
X227 1256 391 390 2 1 1263 QDFFRBN $T=1086860 255480 1 0 $X=1086860 $Y=250060
X228 1265 391 390 2 1 1254 QDFFRBN $T=1105460 225240 1 180 $X=1093680 $Y=224860
X229 1294 391 390 2 1 1277 QDFFRBN $T=1120340 225240 1 180 $X=1108560 $Y=224860
X230 1290 391 403 2 1 1292 QDFFRBN $T=1128400 245400 0 180 $X=1116620 $Y=239980
X231 1287 391 403 2 1 1286 QDFFRBN $T=1128400 245400 1 180 $X=1116620 $Y=245020
X232 1293 391 403 2 1 1296 QDFFRBN $T=1116620 255480 1 0 $X=1116620 $Y=250060
X233 565 55 2 1 56 555 MUX2 $T=343480 255480 0 0 $X=343480 $Y=255100
X234 576 55 2 1 586 59 MUX2 $T=348440 255480 0 0 $X=348440 $Y=255100
X235 585 55 2 1 589 590 MUX2 $T=362080 245400 1 180 $X=357740 $Y=245020
X236 587 55 2 1 599 600 MUX2 $T=362080 245400 0 0 $X=362080 $Y=245020
X237 631 632 639 637 1 634 2 AOI22S $T=414160 235320 0 180 $X=410440 $Y=229900
X238 1160 357 359 1155 1 355 2 AOI22S $T=1029820 255480 0 180 $X=1026100 $Y=250060
X239 354 353 356 1170 1 358 2 AOI22S $T=1026100 255480 0 0 $X=1026100 $Y=255100
X240 365 357 1171 1165 1 363 2 AOI22S $T=1037260 245400 1 180 $X=1033540 $Y=245020
X241 363 357 1177 355 1 364 2 AOI22S $T=1034160 255480 1 0 $X=1034160 $Y=250060
X242 1187 366 1174 364 1 1195 2 AOI22S $T=1037880 245400 1 0 $X=1037880 $Y=239980
X243 1219 366 380 1228 1 1229 2 AOI22S $T=1058960 255480 0 0 $X=1058960 $Y=255100
X244 354 1178 1231 373 1 378 2 AOI22S $T=1063300 255480 0 0 $X=1063300 $Y=255100
X245 626 2 1 73 BUF1 $T=404240 235320 0 180 $X=401760 $Y=229900
X246 94 2 1 648 BUF1 $T=437720 245400 0 0 $X=437720 $Y=245020
X247 102 2 1 52 BUF1 $T=450740 225240 0 180 $X=448260 $Y=219820
X248 107 2 1 671 BUF1 $T=471200 245400 0 0 $X=471200 $Y=245020
X249 118 2 1 677 BUF1 $T=486700 255480 0 180 $X=484220 $Y=250060
X250 156 2 1 741 BUF1 $T=589000 255480 0 180 $X=586520 $Y=250060
X251 189 2 1 802 BUF1 $T=656580 235320 0 180 $X=654100 $Y=229900
X252 192 2 1 810 BUF1 $T=662160 255480 1 180 $X=659680 $Y=255100
X253 198 2 1 811 BUF1 $T=672080 255480 1 0 $X=672080 $Y=250060
X254 302 2 1 102 BUF1 $T=889080 225240 0 180 $X=886600 $Y=219820
X255 405 2 1 54 BUF1 $T=1125300 225240 0 180 $X=1122820 $Y=219820
X256 405 2 1 406 BUF1 $T=1126540 225240 0 0 $X=1126540 $Y=224860
X257 594 1 2 590 BUF1CK $T=365180 245400 1 0 $X=365180 $Y=239980
X258 1078 1 2 314 BUF1CK $T=923800 255480 0 0 $X=923800 $Y=255100
X259 1248 1 2 382 BUF1CK $T=1079420 255480 0 0 $X=1079420 $Y=255100
X260 1263 1 2 1266 BUF1CK $T=1095540 255480 0 0 $X=1095540 $Y=255100
X261 1277 1 2 1280 BUF1CK $T=1104840 235320 0 0 $X=1104840 $Y=234940
X262 184 748 1 2 BUF2 $T=644800 255480 1 0 $X=644800 $Y=250060
X263 625 1 629 630 2 77 ND3 $T=405480 255480 0 0 $X=405480 $Y=255100
X264 207 1 839 837 2 842 ND3 $T=696880 245400 0 0 $X=696880 $Y=245020
X265 841 1 840 824 2 837 ND3 $T=699360 255480 0 180 $X=696880 $Y=250060
X266 826 1 207 840 2 208 ND3 $T=696880 255480 0 0 $X=696880 $Y=255100
X267 826 1 211 849 2 205 ND3 $T=701840 255480 1 0 $X=701840 $Y=250060
X268 859 1 856 218 2 216 ND3 $T=712380 255480 0 0 $X=712380 $Y=255100
X269 851 1 858 866 2 869 ND3 $T=714240 235320 0 0 $X=714240 $Y=234940
X270 1184 1 361 1173 2 354 ND3 $T=1032920 255480 1 180 $X=1030440 $Y=255100
X271 1203 1 361 1202 2 1210 ND3 $T=1044700 255480 0 0 $X=1044700 $Y=255100
X272 1211 1 1207 1198 2 1206 ND3 $T=1049040 245400 0 180 $X=1046560 $Y=239980
X273 1165 1 1187 1211 2 372 ND3 $T=1047180 245400 0 0 $X=1047180 $Y=245020
X274 1232 1 362 1228 2 1231 ND3 $T=1065160 255480 0 180 $X=1062680 $Y=250060
X275 1176 1 1235 1232 2 384 ND3 $T=1067640 255480 1 0 $X=1067640 $Y=250060
X276 383 1 1239 1229 2 1243 ND3 $T=1070120 255480 0 0 $X=1070120 $Y=255100
X277 1264 1 1270 1247 2 1273 ND3 $T=1099880 245400 0 0 $X=1099880 $Y=245020
X278 442 444 8 2 1 ND2S $T=225060 245400 0 180 $X=223200 $Y=239980
X279 444 438 436 2 1 ND2S $T=226920 245400 0 180 $X=225060 $Y=239980
X280 460 461 456 2 1 ND2S $T=247380 225240 1 180 $X=245520 $Y=224860
X281 20 33 450 2 1 ND2S $T=265980 245400 1 180 $X=264120 $Y=245020
X282 530 540 522 2 1 ND2S $T=311860 225240 0 180 $X=310000 $Y=219820
X283 524 522 525 2 1 ND2S $T=310000 225240 0 0 $X=310000 $Y=224860
X284 536 549 545 2 1 ND2S $T=327980 255480 1 180 $X=326120 $Y=255100
X285 548 551 549 2 1 ND2S $T=331080 255480 1 180 $X=329220 $Y=255100
X286 566 570 569 2 1 ND2S $T=340380 255480 1 0 $X=340380 $Y=250060
X287 558 567 571 2 1 ND2S $T=341620 225240 0 0 $X=341620 $Y=224860
X288 535 569 562 2 1 ND2S $T=341620 255480 0 0 $X=341620 $Y=255100
X289 557 579 543 2 1 ND2S $T=347200 225240 0 180 $X=345340 $Y=219820
X290 573 581 567 2 1 ND2S $T=347200 235320 1 180 $X=345340 $Y=234940
X291 578 583 579 2 1 ND2S $T=347820 225240 0 0 $X=347820 $Y=224860
X292 64 574 597 2 1 ND2S $T=360840 235320 0 0 $X=360840 $Y=234940
X293 64 560 598 2 1 ND2S $T=363320 235320 1 0 $X=363320 $Y=229900
X294 596 556 64 2 1 ND2S $T=363320 245400 1 0 $X=363320 $Y=239980
X295 601 559 64 2 1 ND2S $T=366420 245400 0 0 $X=366420 $Y=245020
X296 66 539 64 2 1 ND2S $T=372000 255480 1 180 $X=370140 $Y=255100
X297 76 624 78 2 1 ND2S $T=403620 255480 1 0 $X=403620 $Y=250060
X298 635 633 629 2 1 ND2S $T=411680 255480 0 180 $X=409820 $Y=250060
X299 738 145 737 2 1 ND2S $T=556760 245400 1 180 $X=554900 $Y=245020
X300 831 828 207 2 1 ND2S $T=693780 245400 1 0 $X=693780 $Y=239980
X301 834 832 828 2 1 ND2S $T=693780 255480 1 0 $X=693780 $Y=250060
X302 206 209 205 2 1 ND2S $T=695640 255480 1 180 $X=693780 $Y=255100
X303 836 833 846 2 1 ND2S $T=696880 235320 1 0 $X=696880 $Y=229900
X304 839 838 826 2 1 ND2S $T=698740 245400 1 0 $X=698740 $Y=239980
X305 826 841 845 2 1 ND2S $T=700600 245400 0 0 $X=700600 $Y=245020
X306 827 848 835 2 1 ND2S $T=704320 245400 0 180 $X=702460 $Y=239980
X307 843 846 851 2 1 ND2S $T=704320 235320 1 0 $X=704320 $Y=229900
X308 852 830 854 2 1 ND2S $T=707420 245400 0 0 $X=707420 $Y=245020
X309 852 862 851 2 1 ND2S $T=711140 245400 1 0 $X=711140 $Y=239980
X310 855 867 863 2 1 ND2S $T=716720 245400 1 180 $X=714860 $Y=245020
X311 859 863 217 2 1 ND2S $T=714860 255480 0 0 $X=714860 $Y=255100
X312 868 872 851 2 1 ND2S $T=717960 225240 1 180 $X=716100 $Y=224860
X313 864 875 872 2 1 ND2S $T=722300 225240 0 0 $X=722300 $Y=224860
X314 299 1029 286 2 1 ND2S $T=876680 245400 1 0 $X=876680 $Y=239980
X315 300 1031 1022 2 1 ND2S $T=879780 245400 0 0 $X=879780 $Y=245020
X316 296 1038 1037 2 1 ND2S $T=883500 225240 1 180 $X=881640 $Y=224860
X317 1041 1044 1038 2 1 ND2S $T=884120 235320 0 180 $X=882260 $Y=229900
X318 299 1045 1022 2 1 ND2S $T=885360 255480 0 180 $X=883500 $Y=250060
X319 1042 1046 1044 2 1 ND2S $T=887220 235320 0 180 $X=885360 $Y=229900
X320 297 1049 1037 2 1 ND2S $T=888460 225240 0 0 $X=888460 $Y=224860
X321 296 1050 1043 2 1 ND2S $T=890320 235320 0 180 $X=888460 $Y=229900
X322 300 1047 1034 2 1 ND2S $T=889080 245400 0 0 $X=889080 $Y=245020
X323 1052 1051 296 2 1 ND2S $T=892800 225240 1 180 $X=890940 $Y=224860
X324 300 1041 1052 2 1 ND2S $T=890940 245400 1 0 $X=890940 $Y=239980
X325 1049 1060 1051 2 1 ND2S $T=895900 225240 1 180 $X=894040 $Y=224860
X326 300 1055 1048 2 1 ND2S $T=894040 235320 0 0 $X=894040 $Y=234940
X327 299 1057 1034 2 1 ND2S $T=895900 245400 1 0 $X=895900 $Y=239980
X328 333 1124 332 2 1 ND2S $T=985180 255480 0 180 $X=983320 $Y=250060
X329 337 1127 332 2 1 ND2S $T=991380 255480 0 180 $X=989520 $Y=250060
X330 333 1132 327 2 1 ND2S $T=994480 255480 0 180 $X=992620 $Y=250060
X331 337 1141 327 2 1 ND2S $T=999440 255480 0 180 $X=997580 $Y=250060
X332 333 1143 323 2 1 ND2S $T=1002540 255480 0 180 $X=1000680 $Y=250060
X333 344 1151 349 2 1 ND2S $T=1009980 255480 0 0 $X=1009980 $Y=255100
X334 1165 1155 1176 2 1 ND2S $T=1024240 245400 0 0 $X=1024240 $Y=245020
X335 1160 1180 1168 2 1 ND2S $T=1031060 235320 1 180 $X=1029200 $Y=234940
X336 1179 1162 1186 2 1 ND2S $T=1032920 225240 0 0 $X=1032920 $Y=224860
X337 1188 1190 1180 2 1 ND2S $T=1034780 245400 0 180 $X=1032920 $Y=239980
X338 1160 1184 1194 2 1 ND2S $T=1037880 255480 0 0 $X=1037880 $Y=255100
X339 1197 367 1198 2 1 ND2S $T=1039740 235320 0 0 $X=1039740 $Y=234940
X340 373 1194 1199 2 1 ND2S $T=1045320 255480 1 0 $X=1045320 $Y=250060
X341 1212 1199 374 2 1 ND2S $T=1048420 255480 1 0 $X=1048420 $Y=250060
X342 1190 1220 1216 2 1 ND2S $T=1050900 245400 1 0 $X=1050900 $Y=239980
X343 372 376 1216 2 1 ND2S $T=1050900 255480 1 0 $X=1050900 $Y=250060
X344 371 1203 1222 2 1 ND2S $T=1054000 245400 1 0 $X=1054000 $Y=239980
X345 1219 1210 381 2 1 ND2S $T=1057100 255480 1 0 $X=1057100 $Y=250060
X346 1222 373 1224 2 1 ND2S $T=1065160 235320 0 180 $X=1063300 $Y=229900
X347 1224 1165 365 2 1 ND2S $T=1063300 245400 0 0 $X=1063300 $Y=245020
X348 386 1243 1238 2 1 ND2S $T=1071980 245400 1 180 $X=1070120 $Y=245020
X349 1274 1261 1267 2 1 ND2S $T=1100500 235320 0 0 $X=1100500 $Y=234940
X350 1261 1268 398 2 1 ND2S $T=1102360 235320 1 0 $X=1102360 $Y=229900
X351 1284 1278 1286 2 1 ND2S $T=1107940 255480 1 0 $X=1107940 $Y=250060
X352 399 1282 400 2 1 ND2S $T=1108560 255480 0 0 $X=1108560 $Y=255100
X353 1288 1283 1281 2 1 ND2S $T=1114140 245400 1 0 $X=1114140 $Y=239980
X354 445 8 1 7 443 437 2 MOAI1S $T=227540 245400 1 180 $X=223820 $Y=245020
X355 80 76 1 623 620 621 2 MOAI1S $T=399900 255480 1 180 $X=396180 $Y=255100
X356 638 625 1 82 633 645 2 MOAI1S $T=412300 255480 1 0 $X=412300 $Y=250060
X357 631 636 1 641 628 644 2 MOAI1S $T=412920 235320 0 0 $X=412920 $Y=234940
X358 205 832 1 205 204 203 2 MOAI1S $T=693160 255480 0 180 $X=689440 $Y=250060
X359 827 833 1 827 829 821 2 MOAI1S $T=693780 235320 1 180 $X=690060 $Y=234940
X360 854 867 1 854 862 871 2 MOAI1S $T=716720 245400 1 0 $X=716720 $Y=239980
X361 874 875 1 874 866 877 2 MOAI1S $T=722300 235320 0 0 $X=722300 $Y=234940
X362 1036 287 1 1039 1013 1042 2 MOAI1S $T=880400 245400 1 0 $X=880400 $Y=239980
X363 1050 1059 1 1050 1059 1061 2 MOAI1S $T=895280 235320 1 0 $X=895280 $Y=229900
X364 1055 1057 1 1055 1057 1062 2 MOAI1S $T=897760 235320 0 0 $X=897760 $Y=234940
X365 312 1077 1 312 311 1066 2 MOAI1S $T=923180 255480 0 180 $X=919460 $Y=250060
X366 315 1086 1 315 317 1081 2 MOAI1S $T=931240 255480 0 180 $X=927520 $Y=250060
X367 315 1089 1 315 318 1087 2 MOAI1S $T=935580 255480 0 180 $X=931860 $Y=250060
X368 320 321 1 320 317 1093 2 MOAI1S $T=945500 255480 1 180 $X=941780 $Y=255100
X369 320 322 1 320 311 1099 2 MOAI1S $T=949840 255480 1 180 $X=946120 $Y=255100
X370 1143 1141 1 1143 1141 1145 2 MOAI1S $T=1002540 245400 0 0 $X=1002540 $Y=245020
X371 347 1146 1 347 1146 1149 2 MOAI1S $T=1006260 255480 1 0 $X=1006260 $Y=250060
X372 1151 351 1 1151 351 1146 2 MOAI1S $T=1021140 255480 1 180 $X=1017420 $Y=255100
X373 1155 1160 1 1155 1167 1166 2 MOAI1S $T=1022380 235320 1 0 $X=1022380 $Y=229900
X374 1168 1171 1 1168 1166 1159 2 MOAI1S $T=1028580 225240 1 180 $X=1024860 $Y=224860
X375 1177 1175 1 1173 1172 1153 2 MOAI1S $T=1030440 235320 0 180 $X=1026720 $Y=229900
X376 1187 1185 1 362 1180 1181 2 MOAI1S $T=1034780 235320 0 180 $X=1031060 $Y=229900
X377 1183 1186 1 362 1184 368 2 MOAI1S $T=1034160 255480 0 0 $X=1034160 $Y=255100
X378 1192 1160 1 1189 1188 1185 2 MOAI1S $T=1039120 235320 0 180 $X=1035400 $Y=229900
X379 1169 369 1 1169 1196 1201 2 MOAI1S $T=1039740 235320 1 0 $X=1039740 $Y=229900
X380 353 1202 1 1201 1204 1209 2 MOAI1S $T=1043460 225240 0 0 $X=1043460 $Y=224860
X381 1187 1205 1 1187 1201 1172 2 MOAI1S $T=1047180 235320 1 180 $X=1043460 $Y=234940
X382 371 1192 1 371 1204 1207 2 MOAI1S $T=1050900 235320 0 180 $X=1047180 $Y=229900
X383 1192 1166 1 1214 1189 1218 2 MOAI1S $T=1049660 225240 0 0 $X=1049660 $Y=224860
X384 1192 1220 1 1217 1204 1175 2 MOAI1S $T=1055240 235320 0 180 $X=1051520 $Y=229900
X385 1160 374 1 377 1208 1195 2 MOAI1S $T=1056480 245400 1 180 $X=1052760 $Y=245020
X386 1224 1196 1 1222 371 1221 2 MOAI1S $T=1058960 235320 1 180 $X=1055240 $Y=234940
X387 1222 379 1 1208 1225 1205 2 MOAI1S $T=1056480 245400 1 0 $X=1056480 $Y=239980
X388 1178 1230 1 1227 362 1226 2 MOAI1S $T=1063300 225240 1 180 $X=1059580 $Y=224860
X389 1222 1196 1 1225 369 1230 2 MOAI1S $T=1059580 235320 1 0 $X=1059580 $Y=229900
X390 1176 1196 1 1176 369 1233 2 MOAI1S $T=1063920 225240 0 0 $X=1063920 $Y=224860
X391 1196 1225 1 373 369 1236 2 MOAI1S $T=1065780 235320 1 0 $X=1065780 $Y=229900
X392 1234 385 1 1208 1238 1237 2 MOAI1S $T=1072600 235320 1 180 $X=1068880 $Y=234940
X393 1192 1244 1 1242 1189 1215 2 MOAI1S $T=1075080 225240 1 180 $X=1071360 $Y=224860
X394 365 1234 1 385 1208 1244 2 MOAI1S $T=1073220 235320 0 0 $X=1073220 $Y=234940
X395 1241 1234 1 1241 1208 1249 2 MOAI1S $T=1077560 235320 0 0 $X=1077560 $Y=234940
X396 1161 1247 1 1161 1247 1250 2 MOAI1S $T=1079420 255480 1 0 $X=1079420 $Y=250060
X397 1252 1257 1 1252 1257 1253 2 MOAI1S $T=1091200 235320 1 180 $X=1087480 $Y=234940
X398 1269 1267 1 1264 1251 1256 2 MOAI1S $T=1099260 245400 1 180 $X=1095540 $Y=245020
X399 398 1262 1 1268 1260 1265 2 MOAI1S $T=1101120 235320 0 180 $X=1097400 $Y=229900
X400 1283 1285 1 1283 1285 1291 2 MOAI1S $T=1109180 235320 1 0 $X=1109180 $Y=229900
X401 398 1272 1 402 1289 1293 2 MOAI1S $T=1112900 255480 0 0 $X=1112900 $Y=255100
X402 562 2 563 535 1 NR2 $T=338520 255480 0 180 $X=336660 $Y=250060
X403 543 2 577 557 1 NR2 $T=343480 225240 0 0 $X=343480 $Y=224860
X404 68 2 598 69 1 NR2 $T=375720 235320 1 0 $X=375720 $Y=229900
X405 68 2 593 608 1 NR2 $T=380680 235320 1 0 $X=380680 $Y=229900
X406 68 2 605 609 1 NR2 $T=380680 235320 0 0 $X=380680 $Y=234940
X407 69 2 613 609 1 NR2 $T=380680 245400 1 0 $X=380680 $Y=239980
X408 69 2 606 608 1 NR2 $T=384400 235320 1 0 $X=384400 $Y=229900
X409 68 2 614 71 1 NR2 $T=386260 255480 1 0 $X=386260 $Y=250060
X410 73 2 611 71 1 NR2 $T=389980 255480 1 180 $X=388120 $Y=255100
X411 608 2 604 617 1 NR2 $T=388740 235320 1 0 $X=388740 $Y=229900
X412 72 2 75 609 1 NR2 $T=389980 255480 0 0 $X=389980 $Y=255100
X413 69 2 616 617 1 NR2 $T=390600 235320 1 0 $X=390600 $Y=229900
X414 619 2 615 617 1 NR2 $T=394320 235320 0 180 $X=392460 $Y=229900
X415 626 2 622 609 1 NR2 $T=407340 245400 0 180 $X=405480 $Y=239980
X416 597 2 636 632 1 NR2 $T=406720 235320 0 0 $X=406720 $Y=234940
X417 625 2 635 84 1 NR2 $T=409820 245400 1 180 $X=407960 $Y=245020
X418 635 2 634 638 1 NR2 $T=411060 245400 0 0 $X=411060 $Y=245020
X419 737 2 144 738 1 NR2 $T=554900 255480 1 0 $X=554900 $Y=250060
X420 830 2 206 831 1 NR2 $T=695640 245400 1 180 $X=693780 $Y=245020
X421 209 2 839 210 1 NR2 $T=700600 255480 0 0 $X=700600 $Y=255100
X422 854 2 856 825 1 NR2 $T=709280 245400 0 180 $X=707420 $Y=239980
X423 848 2 858 838 1 NR2 $T=711140 235320 1 180 $X=709280 $Y=234940
X424 214 2 852 859 1 NR2 $T=710520 255480 1 0 $X=710520 $Y=250060
X425 874 2 847 860 1 NR2 $T=721680 235320 1 180 $X=719820 $Y=234940
X426 888 2 889 890 1 NR2 $T=746480 235320 0 0 $X=746480 $Y=234940
X427 888 2 885 233 1 NR2 $T=746480 245400 1 0 $X=746480 $Y=239980
X428 893 2 891 890 1 NR2 $T=748960 245400 1 180 $X=747100 $Y=245020
X429 893 2 895 898 1 NR2 $T=750200 235320 0 0 $X=750200 $Y=234940
X430 894 2 892 233 1 NR2 $T=750200 245400 1 0 $X=750200 $Y=239980
X431 894 2 882 234 1 NR2 $T=750200 245400 0 0 $X=750200 $Y=245020
X432 896 2 900 898 1 NR2 $T=753920 235320 0 0 $X=753920 $Y=234940
X433 888 2 897 902 1 NR2 $T=753920 245400 1 0 $X=753920 $Y=239980
X434 896 2 899 902 1 NR2 $T=753920 245400 0 0 $X=753920 $Y=245020
X435 896 2 903 905 1 NR2 $T=757640 235320 0 180 $X=755780 $Y=229900
X436 898 2 906 236 1 NR2 $T=755780 245400 1 0 $X=755780 $Y=239980
X437 905 2 237 236 1 NR2 $T=755780 255480 0 0 $X=755780 $Y=255100
X438 907 2 904 909 1 NR2 $T=757020 245400 0 0 $X=757020 $Y=245020
X439 888 2 910 898 1 NR2 $T=757640 235320 1 0 $X=757640 $Y=229900
X440 894 2 908 902 1 NR2 $T=760740 245400 0 180 $X=758880 $Y=239980
X441 912 2 238 909 1 NR2 $T=760740 245400 1 180 $X=758880 $Y=245020
X442 912 2 913 234 1 NR2 $T=760120 235320 0 0 $X=760120 $Y=234940
X443 907 2 242 234 1 NR2 $T=762600 245400 1 180 $X=760740 $Y=245020
X444 894 2 914 890 1 NR2 $T=761360 245400 1 0 $X=761360 $Y=239980
X445 907 2 915 233 1 NR2 $T=763220 235320 0 0 $X=763220 $Y=234940
X446 896 2 920 929 1 NR2 $T=773140 235320 1 0 $X=773140 $Y=229900
X447 893 2 919 902 1 NR2 $T=775000 255480 1 0 $X=775000 $Y=250060
X448 929 2 923 236 1 NR2 $T=776860 245400 1 0 $X=776860 $Y=239980
X449 929 2 926 248 1 NR2 $T=776860 245400 0 0 $X=776860 $Y=245020
X450 912 2 930 233 1 NR2 $T=778720 235320 0 0 $X=778720 $Y=234940
X451 907 2 932 890 1 NR2 $T=780580 235320 0 0 $X=780580 $Y=234940
X452 934 2 925 248 1 NR2 $T=782440 245400 1 180 $X=780580 $Y=245020
X453 905 2 935 248 1 NR2 $T=782440 255480 0 180 $X=780580 $Y=250060
X454 936 2 931 909 1 NR2 $T=783680 245400 0 180 $X=781820 $Y=239980
X455 936 2 937 234 1 NR2 $T=784300 235320 1 180 $X=782440 $Y=234940
X456 936 2 928 940 1 NR2 $T=784300 245400 0 0 $X=784300 $Y=245020
X457 912 2 939 940 1 NR2 $T=784300 255480 1 0 $X=784300 $Y=250060
X458 912 2 943 890 1 NR2 $T=785540 235320 0 0 $X=785540 $Y=234940
X459 936 2 933 942 1 NR2 $T=786780 255480 1 0 $X=786780 $Y=250060
X460 942 2 922 945 1 NR2 $T=788640 255480 1 0 $X=788640 $Y=250060
X461 257 2 918 253 1 NR2 $T=792360 255480 0 0 $X=792360 $Y=255100
X462 934 2 947 236 1 NR2 $T=792980 245400 0 0 $X=792980 $Y=245020
X463 909 2 946 945 1 NR2 $T=792980 255480 1 0 $X=792980 $Y=250060
X464 894 2 950 898 1 NR2 $T=795460 245400 1 0 $X=795460 $Y=239980
X465 893 2 261 905 1 NR2 $T=796080 255480 0 0 $X=796080 $Y=255100
X466 955 2 949 248 1 NR2 $T=799800 245400 1 180 $X=797940 $Y=245020
X467 896 2 953 934 1 NR2 $T=798560 245400 1 0 $X=798560 $Y=239980
X468 234 2 957 945 1 NR2 $T=801660 235320 0 0 $X=801660 $Y=234940
X469 955 2 958 236 1 NR2 $T=801660 245400 1 0 $X=801660 $Y=239980
X470 936 2 960 233 1 NR2 $T=805380 235320 0 0 $X=805380 $Y=234940
X471 907 2 961 902 1 NR2 $T=808480 245400 1 0 $X=808480 $Y=239980
X472 963 2 962 905 1 NR2 $T=812820 245400 0 180 $X=810960 $Y=239980
X473 963 2 965 934 1 NR2 $T=812820 245400 1 0 $X=812820 $Y=239980
X474 966 2 964 929 1 NR2 $T=814680 245400 1 180 $X=812820 $Y=245020
X475 966 2 970 934 1 NR2 $T=817160 255480 0 180 $X=815300 $Y=250060
X476 966 2 967 955 1 NR2 $T=815920 245400 1 0 $X=815920 $Y=239980
X477 896 2 973 955 1 NR2 $T=815920 245400 0 0 $X=815920 $Y=245020
X478 890 2 976 945 1 NR2 $T=819640 245400 1 0 $X=819640 $Y=239980
X479 233 2 974 945 1 NR2 $T=819640 255480 1 0 $X=819640 $Y=250060
X480 902 2 272 236 1 NR2 $T=823360 255480 0 180 $X=821500 $Y=250060
X481 936 2 980 274 1 NR2 $T=826460 255480 0 180 $X=824600 $Y=250060
X482 977 2 978 905 1 NR2 $T=828320 245400 0 180 $X=826460 $Y=239980
X483 907 2 979 898 1 NR2 $T=826460 245400 0 0 $X=826460 $Y=245020
X484 963 2 988 929 1 NR2 $T=832040 235320 0 0 $X=832040 $Y=234940
X485 992 2 990 985 1 NR2 $T=837000 245400 1 180 $X=835140 $Y=245020
X486 977 2 989 929 1 NR2 $T=835760 235320 0 0 $X=835760 $Y=234940
X487 912 2 983 278 1 NR2 $T=835760 245400 1 0 $X=835760 $Y=239980
X488 987 2 991 985 1 NR2 $T=838860 235320 0 0 $X=838860 $Y=234940
X489 963 2 997 955 1 NR2 $T=840720 235320 0 0 $X=840720 $Y=234940
X490 996 2 285 998 1 NR2 $T=841960 255480 1 0 $X=841960 $Y=250060
X491 985 2 999 945 1 NR2 $T=843200 235320 0 0 $X=843200 $Y=234940
X492 977 2 1002 934 1 NR2 $T=847540 245400 0 180 $X=845680 $Y=239980
X493 977 2 1003 1004 1 NR2 $T=847540 235320 0 0 $X=847540 $Y=234940
X494 996 2 1005 1007 1 NR2 $T=851880 245400 1 0 $X=851880 $Y=239980
X495 278 2 1010 287 1 NR2 $T=856840 245400 0 180 $X=854980 $Y=239980
X496 996 2 1014 1013 1 NR2 $T=856840 235320 1 0 $X=856840 $Y=229900
X497 996 2 1012 955 1 NR2 $T=856840 245400 1 0 $X=856840 $Y=239980
X498 987 2 1015 278 1 NR2 $T=860560 235320 0 180 $X=858700 $Y=229900
X499 987 2 1016 1013 1 NR2 $T=863040 245400 1 180 $X=861180 $Y=245020
X500 1013 2 1020 287 1 NR2 $T=861800 245400 1 0 $X=861800 $Y=239980
X501 992 2 1011 998 1 NR2 $T=864280 235320 1 0 $X=864280 $Y=229900
X502 998 2 1019 287 1 NR2 $T=866140 255480 1 0 $X=866140 $Y=250060
X503 992 2 1023 1013 1 NR2 $T=867380 235320 1 0 $X=867380 $Y=229900
X504 992 2 1028 1004 1 NR2 $T=869240 235320 1 0 $X=869240 $Y=229900
X505 987 2 1026 1007 1 NR2 $T=869240 245400 1 0 $X=869240 $Y=239980
X506 992 2 1024 1007 1 NR2 $T=869240 255480 1 0 $X=869240 $Y=250060
X507 1031 2 1027 1029 1 NR2 $T=874820 245400 0 0 $X=874820 $Y=245020
X508 987 2 1032 998 1 NR2 $T=876680 235320 1 0 $X=876680 $Y=229900
X509 1004 2 1043 1041 1 NR2 $T=881640 235320 0 0 $X=881640 $Y=234940
X510 1047 2 1035 1045 1 NR2 $T=887220 245400 1 180 $X=885360 $Y=245020
X511 1055 2 1054 1057 1 NR2 $T=894040 245400 1 0 $X=894040 $Y=239980
X512 1124 2 1123 335 1 NR2 $T=988280 255480 0 180 $X=986420 $Y=250060
X513 1132 2 1131 1127 1 NR2 $T=993860 245400 1 180 $X=992000 $Y=245020
X514 338 2 1125 339 1 NR2 $T=992000 255480 0 0 $X=992000 $Y=255100
X515 341 2 1128 340 1 NR2 $T=996340 255480 1 180 $X=994480 $Y=255100
X516 342 2 1129 340 1 NR2 $T=1000680 255480 1 180 $X=998820 $Y=255100
X517 1143 2 1142 1141 1 NR2 $T=1002540 245400 1 180 $X=1000680 $Y=245020
X518 342 2 1139 339 1 NR2 $T=1002540 255480 1 180 $X=1000680 $Y=255100
X519 346 2 1144 340 1 NR2 $T=1006260 255480 0 180 $X=1004400 $Y=250060
X520 1157 2 1164 1163 1 NR2 $T=1021760 235320 0 0 $X=1021760 $Y=234940
X521 1169 2 1163 1167 1 NR2 $T=1026100 235320 0 0 $X=1026100 $Y=234940
X522 1189 2 1183 1188 1 NR2 $T=1036640 235320 1 180 $X=1034780 $Y=234940
X523 370 2 363 371 1 NR2 $T=1041600 255480 0 0 $X=1041600 $Y=255100
X524 372 2 1219 371 1 NR2 $T=1052140 255480 0 0 $X=1052140 $Y=255100
X525 1157 2 1214 1221 1 NR2 $T=1054000 225240 0 0 $X=1054000 $Y=224860
X526 378 2 1186 374 1 NR2 $T=1055860 255480 0 180 $X=1054000 $Y=250060
X527 1224 2 1157 369 1 NR2 $T=1059580 235320 0 0 $X=1059580 $Y=234940
X528 1222 2 377 1224 1 NR2 $T=1060820 245400 1 0 $X=1060820 $Y=239980
X529 1224 2 1225 365 1 NR2 $T=1062680 235320 0 0 $X=1062680 $Y=234940
X530 1161 2 1178 382 1 NR2 $T=1065160 255480 1 0 $X=1065160 $Y=250060
X531 1233 2 1227 1237 1 NR2 $T=1068260 225240 0 0 $X=1068260 $Y=224860
X532 1235 2 353 382 1 NR2 $T=1070120 245400 1 180 $X=1068260 $Y=245020
X533 1238 2 1217 1240 1 NR2 $T=1070120 235320 1 0 $X=1070120 $Y=229900
X534 1234 2 1240 1196 1 NR2 $T=1073840 235320 0 180 $X=1071980 $Y=229900
X535 1235 2 386 389 1 NR2 $T=1076940 255480 1 0 $X=1076940 $Y=250060
X536 1161 2 388 389 1 NR2 $T=1076940 255480 0 0 $X=1076940 $Y=255100
X537 1249 2 1242 1236 1 NR2 $T=1081900 235320 0 0 $X=1081900 $Y=234940
X538 1251 2 1255 1253 1 NR2 $T=1084380 235320 0 0 $X=1084380 $Y=234940
X539 1251 2 1258 1250 1 NR2 $T=1086240 245400 1 180 $X=1084380 $Y=245020
X540 1260 2 1257 1261 1 NR2 $T=1091200 235320 1 0 $X=1091200 $Y=229900
X541 1259 2 1262 1261 1 NR2 $T=1094920 235320 0 0 $X=1094920 $Y=234940
X542 1274 2 1269 393 1 NR2 $T=1098640 235320 1 180 $X=1096780 $Y=234940
X543 1283 2 1274 1285 1 NR2 $T=1107320 235320 0 0 $X=1107320 $Y=234940
X544 401 2 399 1289 1 NR2 $T=1111040 255480 0 0 $X=1111040 $Y=255100
X545 1291 2 1294 393 1 NR2 $T=1117860 235320 0 180 $X=1116000 $Y=229900
X546 1295 2 1272 401 1 NR2 $T=1119100 255480 1 180 $X=1117240 $Y=255100
X547 484 475 2 1 502 OR2 $T=275900 235320 1 0 $X=275900 $Y=229900
X548 524 525 2 1 530 OR2 $T=309380 235320 1 0 $X=309380 $Y=229900
X549 536 545 2 1 548 OR2 $T=325500 255480 1 0 $X=325500 $Y=250060
X550 558 571 2 1 573 OR2 $T=341620 235320 1 0 $X=341620 $Y=229900
X551 82 630 2 1 632 OR2 $T=406100 255480 1 0 $X=406100 $Y=250060
X552 91 87 2 1 646 OR2 $T=430900 255480 0 180 $X=428420 $Y=250060
X553 647 654 2 1 657 OR2 $T=444540 225240 0 0 $X=444540 $Y=224860
X554 665 678 2 1 692 OR2 $T=487320 225240 0 0 $X=487320 $Y=224860
X555 698 693 2 1 176 OR2 $T=623720 245400 0 0 $X=623720 $Y=245020
X556 1215 1209 2 1 1200 OR2 $T=1049040 225240 0 180 $X=1046560 $Y=219820
X557 1226 1218 2 1 1193 OR2 $T=1059580 225240 1 180 $X=1057100 $Y=224860
X558 1267 1271 2 1 1264 OR2 $T=1102360 245400 0 180 $X=1099880 $Y=239980
X559 503 45 1 2 532 AN2 $T=302560 225240 1 0 $X=302560 $Y=219820
X560 500 45 1 2 516 AN2 $T=302560 225240 0 0 $X=302560 $Y=224860
X561 508 45 1 2 526 AN2 $T=305660 235320 1 0 $X=305660 $Y=229900
X562 511 45 1 2 529 AN2 $T=307520 245400 1 0 $X=307520 $Y=239980
X563 507 45 1 2 531 AN2 $T=310000 235320 0 0 $X=310000 $Y=234940
X564 1272 2 395 1275 1273 1 NR3 $T=1101120 255480 0 0 $X=1101120 $Y=255100
X565 1262 2 396 1276 1270 1 NR3 $T=1102980 255480 1 0 $X=1102980 $Y=250060
X566 517 48 1 533 2 OR2B1S $T=313720 235320 0 0 $X=313720 $Y=234940
X567 761 156 1 752 2 OR2B1S $T=583420 255480 0 180 $X=580320 $Y=250060
X568 761 811 1 814 2 OR2B1S $T=670220 245400 0 0 $X=670220 $Y=245020
X569 400 399 1 397 2 OR2B1S $T=1108560 255480 1 180 $X=1105460 $Y=255100
X570 755 154 756 1 2 ND2 $T=575980 255480 0 0 $X=575980 $Y=255100
X571 764 159 762 1 2 ND2 $T=589000 255480 1 0 $X=589000 $Y=250060
X572 398 1283 1288 1281 2 1 1290 OA112 $T=1110420 235320 0 0 $X=1110420 $Y=234940
X573 398 1278 1284 1286 2 1 1279 OA112 $T=1110420 255480 1 0 $X=1110420 $Y=250060
X574 1180 1176 1 1174 1170 1164 2 OAI112HS $T=1031680 245400 0 180 $X=1027340 $Y=239980
X575 756 2 755 1 155 NR2P $T=579080 255480 0 0 $X=579080 $Y=255100
X576 762 2 764 1 157 NR2P $T=589620 255480 1 180 $X=585900 $Y=255100
X577 843 842 847 2 827 1 213 AN4B1S $T=701840 235320 0 0 $X=701840 $Y=234940
X578 1162 1159 353 2 1157 1 1154 AN4B1S $T=1024240 225240 1 180 $X=1019900 $Y=224860
X579 492 2 485 478 474 1 499 FA1S $T=268460 225240 1 0 $X=268460 $Y=219820
X580 496 2 488 477 40 1 504 FA1S $T=275280 245400 1 0 $X=275280 $Y=239980
X581 498 2 39 476 494 1 42 FA1S $T=276520 255480 0 0 $X=276520 $Y=255100
X582 500 2 490 497 499 1 510 FA1S $T=278380 225240 0 0 $X=278380 $Y=224860
X583 497 2 467 479 495 1 505 FA1S $T=279000 235320 0 0 $X=279000 $Y=234940
X584 501 2 491 462 498 1 506 FA1S $T=279620 245400 0 0 $X=279620 $Y=245020
X585 503 2 482 493 492 1 514 FA1S $T=284580 225240 1 0 $X=284580 $Y=219820
X586 507 2 496 505 501 1 515 FA1S $T=289540 245400 1 0 $X=289540 $Y=239980
X587 508 2 487 489 486 1 518 FA1S $T=290160 235320 1 0 $X=290160 $Y=229900
X588 509 2 465 41 43 1 44 FA1S $T=291400 255480 0 0 $X=291400 $Y=255100
X589 511 2 504 506 509 1 520 FA1S $T=293880 245400 0 0 $X=293880 $Y=245020
X590 535 2 529 538 537 1 545 FA1S $T=311240 245400 0 0 $X=311240 $Y=245020
X591 537 2 542 539 527 1 528 FA1S $T=324260 255480 0 180 $X=312480 $Y=250060
X592 536 2 47 528 49 1 50 FA1S $T=312480 255480 0 0 $X=312480 $Y=255100
X593 524 2 532 534 544 1 543 FA1S $T=313100 225240 0 0 $X=313100 $Y=224860
X594 541 2 574 572 523 1 534 FA1S $T=329840 235320 1 180 $X=318060 $Y=234940
X595 553 2 564 559 519 1 538 FA1S $T=337280 245400 1 180 $X=325500 $Y=245020
X596 544 2 560 568 521 1 546 FA1S $T=339140 225240 1 180 $X=327360 $Y=224860
X597 554 2 561 556 513 1 547 FA1S $T=339140 235320 0 180 $X=327360 $Y=229900
X598 557 2 516 546 554 1 571 FA1S $T=332320 225240 1 0 $X=332320 $Y=219820
X599 558 2 531 547 553 1 562 FA1S $T=332940 245400 1 0 $X=332940 $Y=239980
X600 596 2 605 604 603 1 588 FA1S $T=378200 235320 1 180 $X=366420 $Y=234940
X601 595 2 612 615 606 1 591 FA1S $T=383780 225240 1 180 $X=372000 $Y=224860
X602 601 2 614 607 610 1 582 FA1S $T=385640 255480 0 180 $X=373860 $Y=250060
X603 607 2 70 613 611 1 67 FA1S $T=385640 255480 1 180 $X=373860 $Y=255100
X604 603 2 74 616 622 1 610 FA1S $T=399900 235320 1 180 $X=388120 $Y=234940
X605 652 2 649 93 98 1 659 FA1S $T=436480 255480 1 0 $X=436480 $Y=250060
X606 700 2 682 666 694 1 707 FA1S $T=494760 245400 0 0 $X=494760 $Y=245020
X607 705 2 688 695 702 1 710 FA1S $T=500340 225240 0 0 $X=500340 $Y=224860
X608 712 2 652 676 129 1 131 FA1S $T=512740 255480 1 0 $X=512740 $Y=250060
X609 715 2 706 672 130 1 718 FA1S $T=515220 235320 1 0 $X=515220 $Y=229900
X610 719 2 135 707 133 1 137 FA1S $T=525140 255480 0 0 $X=525140 $Y=255100
X611 721 2 719 708 717 1 726 FA1S $T=525760 255480 1 0 $X=525760 $Y=250060
X612 725 2 729 722 732 1 736 FA1S $T=532580 225240 0 0 $X=532580 $Y=224860
X613 727 2 723 720 728 1 733 FA1S $T=535680 235320 0 0 $X=535680 $Y=234940
X614 142 2 735 731 727 1 738 FA1S $T=546840 245400 1 0 $X=546840 $Y=239980
X615 739 2 683 150 146 1 732 FA1S $T=562340 235320 1 180 $X=550560 $Y=234940
X616 751 2 757 758 746 1 747 FA1S $T=576600 235320 1 180 $X=564820 $Y=234940
X617 766 2 771 710 161 1 740 FA1S $T=597060 225240 1 180 $X=585280 $Y=224860
X618 769 2 768 167 703 1 782 FA1S $T=590860 245400 1 0 $X=590860 $Y=239980
X619 774 2 778 705 770 1 781 FA1S $T=597060 235320 1 0 $X=597060 $Y=229900
X620 775 2 780 769 774 1 765 FA1S $T=608840 235320 1 180 $X=597060 $Y=234940
X621 779 2 766 782 781 1 759 FA1S $T=611940 225240 1 180 $X=600160 $Y=224860
X622 783 2 791 174 716 1 780 FA1S $T=623100 235320 1 180 $X=611320 $Y=234940
X623 784 2 792 794 179 1 790 FA1S $T=634260 245400 0 180 $X=622480 $Y=239980
X624 793 2 177 772 798 1 796 FA1S $T=627440 255480 1 0 $X=627440 $Y=250060
X625 799 2 803 800 182 1 757 FA1S $T=646660 235320 1 180 $X=634880 $Y=234940
X626 188 2 809 191 808 1 797 FA1S $T=656580 255480 1 180 $X=644800 $Y=255100
X627 228 2 883 884 878 1 224 FA1S $T=744000 255480 0 180 $X=732220 $Y=250060
X628 229 2 880 886 881 1 225 FA1S $T=745240 225240 0 180 $X=733460 $Y=219820
X629 230 2 885 891 882 1 878 FA1S $T=746480 245400 1 180 $X=734700 $Y=245020
X630 231 2 901 887 232 1 226 FA1S $T=749580 255480 1 180 $X=737800 $Y=255100
X631 887 2 889 900 892 1 880 FA1S $T=752060 235320 0 180 $X=740280 $Y=229900
X632 235 2 899 906 904 1 883 FA1S $T=758260 255480 0 180 $X=746480 $Y=250060
X633 886 2 903 895 897 1 911 FA1S $T=747720 225240 1 0 $X=747720 $Y=219820
X634 244 2 919 917 918 1 240 FA1S $T=771280 255480 1 180 $X=759500 $Y=255100
X635 245 2 921 916 911 1 241 FA1S $T=771900 235320 0 180 $X=760120 $Y=229900
X636 916 2 920 910 908 1 924 FA1S $T=762600 225240 1 0 $X=762600 $Y=219820
X637 901 2 926 928 922 1 243 FA1S $T=775620 245400 1 180 $X=763840 $Y=245020
X638 917 2 914 923 925 1 246 FA1S $T=764460 245400 1 0 $X=764460 $Y=239980
X639 881 2 913 915 931 1 247 FA1S $T=765700 235320 0 0 $X=765700 $Y=234940
X640 250 2 939 935 933 1 884 FA1S $T=784920 255480 1 180 $X=773140 $Y=255100
X641 921 2 932 930 937 1 927 FA1S $T=787400 225240 1 180 $X=775620 $Y=224860
X642 251 2 938 924 927 1 941 FA1S $T=776860 225240 1 0 $X=776860 $Y=219820
X643 255 2 947 949 946 1 938 FA1S $T=795460 245400 0 180 $X=783680 $Y=239980
X644 260 2 948 956 951 1 944 FA1S $T=801660 225240 1 180 $X=789880 $Y=224860
X645 948 2 943 950 953 1 954 FA1S $T=789880 235320 0 0 $X=789880 $Y=234940
X646 259 2 941 944 959 1 264 FA1S $T=791740 225240 1 0 $X=791740 $Y=219820
X647 263 2 952 954 968 1 267 FA1S $T=797940 255480 0 0 $X=797940 $Y=255100
X648 956 2 962 964 961 1 952 FA1S $T=812820 245400 1 180 $X=801040 $Y=245020
X649 951 2 960 958 957 1 972 FA1S $T=804140 225240 0 0 $X=804140 $Y=224860
X650 959 2 972 975 969 1 266 FA1S $T=818400 225240 0 180 $X=806620 $Y=219820
X651 971 2 965 967 976 1 982 FA1S $T=812200 235320 0 0 $X=812200 $Y=234940
X652 271 2 973 970 974 1 275 FA1S $T=814680 255480 0 0 $X=814680 $Y=255100
X653 969 2 981 269 971 1 984 FA1S $T=818400 225240 0 0 $X=818400 $Y=224860
X654 280 2 993 984 986 1 273 FA1S $T=836380 225240 0 180 $X=824600 $Y=219820
X655 975 2 988 277 978 1 993 FA1S $T=826460 235320 1 0 $X=826460 $Y=229900
X656 968 2 979 990 980 1 282 FA1S $T=827700 255480 1 0 $X=827700 $Y=250060
X657 281 2 982 279 284 1 995 FA1S $T=830180 255480 0 0 $X=830180 $Y=255100
X658 981 2 983 991 989 1 1000 FA1S $T=833900 225240 0 0 $X=833900 $Y=224860
X659 986 2 1000 1008 1001 1 994 FA1S $T=853120 225240 0 180 $X=841340 $Y=219820
X660 1001 2 1002 997 999 1 1006 FA1S $T=841340 235320 1 0 $X=841340 $Y=229900
X661 288 2 995 994 1009 1 291 FA1S $T=844440 255480 0 0 $X=844440 $Y=255100
X662 290 2 1005 1003 1010 1 294 FA1S $T=849400 255480 1 0 $X=849400 $Y=250060
X663 1009 2 1006 1021 1018 1 289 FA1S $T=863660 225240 1 180 $X=851880 $Y=224860
X664 1008 2 1014 1011 1015 1 1021 FA1S $T=856220 225240 1 0 $X=856220 $Y=219820
X665 293 2 1016 1012 1019 1 1025 FA1S $T=858080 255480 0 0 $X=858080 $Y=255100
X666 1018 2 1027 1023 1032 1 295 FA1S $T=879780 225240 1 180 $X=868000 $Y=224860
X667 298 2 1030 1035 1024 1 1040 FA1S $T=871100 255480 1 0 $X=871100 $Y=250060
X668 301 2 1033 1040 1025 1 303 FA1S $T=881640 255480 0 0 $X=881640 $Y=255100
X669 304 2 1017 1053 1054 1 1063 FA1S $T=892180 245400 0 0 $X=892180 $Y=245020
X670 305 2 1058 1056 1064 1 307 FA1S $T=895900 255480 0 0 $X=895900 $Y=255100
X671 309 2 313 1080 1076 1 1065 FA1S $T=924420 245400 1 180 $X=912640 $Y=245020
X672 1076 2 1077 1083 1079 1 1070 FA1S $T=927520 245400 0 180 $X=915740 $Y=239980
X673 1079 2 1086 1084 1082 1 1068 FA1S $T=930620 235320 0 180 $X=918840 $Y=229900
X674 1082 2 1078 1092 1085 1 1074 FA1S $T=933100 225240 1 180 $X=921320 $Y=224860
X675 1085 2 319 1089 1094 1 1088 FA1S $T=943020 235320 0 180 $X=931240 $Y=229900
X676 325 2 1107 324 1106 1 1108 FA1S $T=952320 255480 0 0 $X=952320 $Y=255100
X677 1107 2 326 328 1112 1 1116 FA1S $T=964720 255480 0 0 $X=964720 $Y=255100
X678 1106 2 1113 1116 1115 1 1110 FA1S $T=980220 235320 1 180 $X=968440 $Y=234940
X679 1113 2 1119 1118 1114 1 1109 FA1S $T=980220 245400 0 180 $X=968440 $Y=239980
X680 1112 2 330 329 331 1 1118 FA1S $T=968440 255480 1 0 $X=968440 $Y=250060
X681 1115 2 1121 1109 1117 1 1111 FA1S $T=982080 235320 0 180 $X=970300 $Y=229900
X682 334 2 1123 1128 1125 1 1114 FA1S $T=990140 255480 1 180 $X=978360 $Y=255100
X683 1119 2 1126 1131 1129 1 1120 FA1S $T=994480 245400 0 180 $X=982700 $Y=239980
X684 1117 2 1135 1134 1130 1 1122 FA1S $T=995720 225240 1 180 $X=983940 $Y=224860
X685 1121 2 1133 1120 336 1 1134 FA1S $T=983940 235320 1 0 $X=983940 $Y=229900
X686 1133 2 1144 1139 343 1 1138 FA1S $T=1009360 245400 0 180 $X=997580 $Y=239980
X687 1130 2 1138 1136 1142 1 1140 FA1S $T=998820 235320 1 0 $X=998820 $Y=229900
X688 16 17 457 2 1 XNR2HS $T=241180 245400 0 0 $X=241180 $Y=245020
X689 16 18 458 2 1 XNR2HS $T=249240 255480 1 180 $X=243660 $Y=255100
X690 452 450 20 2 1 XNR2HS $T=245520 245400 1 0 $X=245520 $Y=239980
X691 463 18 466 2 1 XNR2HS $T=248620 225240 0 0 $X=248620 $Y=224860
X692 463 24 468 2 1 XNR2HS $T=250480 235320 0 0 $X=250480 $Y=234940
X693 463 26 470 2 1 XNR2HS $T=254820 245400 1 0 $X=254820 $Y=239980
X694 463 17 471 2 1 XNR2HS $T=255440 225240 0 0 $X=255440 $Y=224860
X695 25 27 472 2 1 XNR2HS $T=255440 255480 0 0 $X=255440 $Y=255100
X696 551 53 565 2 1 XNR2HS $T=336040 255480 0 0 $X=336040 $Y=255100
X697 581 584 585 2 1 XNR2HS $T=349060 245400 1 0 $X=349060 $Y=239980
X698 92 90 88 2 1 XNR2HS $T=434620 255480 1 180 $X=429040 $Y=255100
X699 87 91 649 2 1 XNR2HS $T=432140 245400 0 0 $X=432140 $Y=245020
X700 92 648 650 2 1 XNR2HS $T=433380 235320 0 0 $X=433380 $Y=234940
X701 95 648 653 2 1 XNR2HS $T=437720 245400 1 0 $X=437720 $Y=239980
X702 103 648 97 2 1 XNR2HS $T=450740 245400 1 180 $X=445160 $Y=245020
X703 654 647 660 2 1 XNR2HS $T=448260 225240 0 0 $X=448260 $Y=224860
X704 92 104 661 2 1 XNR2HS $T=448880 235320 0 0 $X=448880 $Y=234940
X705 106 104 662 2 1 XNR2HS $T=453840 245400 0 0 $X=453840 $Y=245020
X706 95 104 663 2 1 XNR2HS $T=456320 235320 0 0 $X=456320 $Y=234940
X707 111 112 673 2 1 XNR2HS $T=464380 255480 0 0 $X=464380 $Y=255100
X708 103 104 668 2 1 XNR2HS $T=465000 245400 1 0 $X=465000 $Y=239980
X709 95 112 674 2 1 XNR2HS $T=465000 245400 0 0 $X=465000 $Y=245020
X710 103 116 684 2 1 XNR2HS $T=475540 245400 1 0 $X=475540 $Y=239980
X711 106 116 686 2 1 XNR2HS $T=482980 245400 0 0 $X=482980 $Y=245020
X712 92 116 690 2 1 XNR2HS $T=482980 255480 0 0 $X=482980 $Y=255100
X713 678 665 695 2 1 XNR2HS $T=491040 225240 0 0 $X=491040 $Y=224860
X714 125 127 704 2 1 XNR2HS $T=499720 255480 0 0 $X=499720 $Y=255100
X715 147 741 744 2 1 XNR2HS $T=558000 255480 1 0 $X=558000 $Y=250060
X716 151 741 745 2 1 XNR2HS $T=574120 255480 0 180 $X=568540 $Y=250060
X717 158 741 749 2 1 XNR2HS $T=589000 245400 1 180 $X=583420 $Y=245020
X718 693 698 792 2 1 XNR2HS $T=626200 235320 0 0 $X=626200 $Y=234940
X719 180 156 760 2 1 XNR2HS $T=641080 245400 0 180 $X=635500 $Y=239980
X720 181 156 801 2 1 XNR2HS $T=639220 255480 1 0 $X=639220 $Y=250060
X721 761 810 807 2 1 XNR2HS $T=659060 225240 1 180 $X=653480 $Y=224860
X722 158 810 804 2 1 XNR2HS $T=659060 235320 1 180 $X=653480 $Y=234940
X723 180 810 806 2 1 XNR2HS $T=659060 245400 1 180 $X=653480 $Y=245020
X724 181 810 190 2 1 XNR2HS $T=660920 255480 0 180 $X=655340 $Y=250060
X725 147 810 805 2 1 XNR2HS $T=658440 235320 1 0 $X=658440 $Y=229900
X726 147 811 812 2 1 XNR2HS $T=660300 235320 0 0 $X=660300 $Y=234940
X727 158 811 813 2 1 XNR2HS $T=660920 255480 1 0 $X=660920 $Y=250060
X728 761 811 815 2 1 XNR2HS $T=667120 235320 0 0 $X=667120 $Y=234940
X729 180 198 197 2 1 XNR2HS $T=670840 255480 0 0 $X=670840 $Y=255100
X730 76 82 78 1 2 623 OA12 $T=403000 255480 0 180 $X=399280 $Y=250060
X731 84 631 634 1 2 641 OA12 $T=411060 245400 1 0 $X=411060 $Y=239980
X732 1048 1043 299 1 2 1036 OA12 $T=887840 245400 0 180 $X=884120 $Y=239980
X733 1049 1051 1050 1 2 1056 OA12 $T=890940 235320 1 0 $X=890940 $Y=229900
X734 21 1 457 19 462 458 2 OAI22S $T=251100 245400 1 180 $X=247380 $Y=245020
X735 21 1 458 19 465 23 2 OAI22S $T=254820 255480 1 180 $X=251100 $Y=255100
X736 22 1 21 19 467 457 2 OAI22S $T=255440 245400 1 180 $X=251720 $Y=245020
X737 460 1 466 461 479 468 2 OAI22S $T=260400 235320 0 0 $X=260400 $Y=234940
X738 480 1 470 31 476 472 2 OAI22S $T=264740 255480 0 180 $X=261020 $Y=250060
X739 32 1 472 31 30 29 2 OAI22S $T=264740 255480 1 180 $X=261020 $Y=255100
X740 480 1 468 461 477 470 2 OAI22S $T=265360 245400 0 180 $X=261640 $Y=239980
X741 460 1 471 461 478 466 2 OAI22S $T=265980 225240 1 180 $X=262260 $Y=224860
X742 473 1 481 484 485 483 2 OAI22S $T=266600 245400 1 0 $X=266600 $Y=239980
X743 28 1 460 461 482 471 2 OAI22S $T=270940 225240 1 180 $X=267220 $Y=224860
X744 464 1 481 484 487 469 2 OAI22S $T=267220 235320 0 0 $X=267220 $Y=234940
X745 35 1 481 33 488 36 2 OAI22S $T=268460 255480 1 0 $X=268460 $Y=250060
X746 483 1 481 484 491 35 2 OAI22S $T=269700 245400 0 0 $X=269700 $Y=245020
X747 475 1 481 484 489 464 2 OAI22S $T=274660 235320 0 180 $X=270940 $Y=229900
X748 469 1 481 484 490 473 2 OAI22S $T=274660 245400 0 180 $X=270940 $Y=239980
X749 36 1 20 33 37 38 2 OAI22S $T=271560 255480 0 0 $X=271560 $Y=255100
X750 96 1 650 653 654 99 2 OAI22S $T=439580 235320 0 0 $X=439580 $Y=234940
X751 96 1 653 97 655 100 2 OAI22S $T=440820 245400 0 0 $X=440820 $Y=245020
X752 110 1 662 109 664 107 2 OAI22S $T=464380 245400 1 180 $X=460660 $Y=245020
X753 110 1 668 662 669 671 2 OAI22S $T=462520 235320 0 0 $X=462520 $Y=234940
X754 110 1 663 668 675 671 2 OAI22S $T=466860 235320 0 0 $X=466860 $Y=234940
X755 110 1 661 663 678 671 2 OAI22S $T=471200 235320 0 0 $X=471200 $Y=234940
X756 677 1 673 113 667 680 2 OAI22S $T=471200 255480 1 0 $X=471200 $Y=250060
X757 677 1 114 115 681 680 2 OAI22S $T=474300 245400 0 0 $X=474300 $Y=245020
X758 677 1 115 673 682 680 2 OAI22S $T=475540 255480 1 0 $X=475540 $Y=250060
X759 677 1 686 114 685 680 2 OAI22S $T=482360 245400 1 180 $X=478640 $Y=245020
X760 118 1 684 686 688 687 2 OAI22S $T=481740 245400 1 0 $X=481740 $Y=239980
X761 118 1 674 684 691 687 2 OAI22S $T=486080 245400 1 0 $X=486080 $Y=239980
X762 118 1 690 674 693 687 2 OAI22S $T=492900 245400 1 180 $X=489180 $Y=245020
X763 120 1 121 122 694 123 2 OAI22S $T=491660 255480 1 0 $X=491660 $Y=250060
X764 120 1 124 122 697 121 2 OAI22S $T=499720 255480 0 180 $X=496000 $Y=250060
X765 120 1 126 122 702 704 2 OAI22S $T=499720 255480 1 0 $X=499720 $Y=250060
X766 120 1 704 122 706 124 2 OAI22S $T=504060 255480 1 0 $X=504060 $Y=250060
X767 120 1 128 122 709 126 2 OAI22S $T=508400 255480 1 0 $X=508400 $Y=250060
X768 748 1 744 148 714 745 2 OAI22S $T=566680 245400 1 180 $X=562960 $Y=245020
X769 748 1 749 148 730 744 2 OAI22S $T=571020 245400 1 180 $X=567300 $Y=245020
X770 753 1 148 752 724 748 2 OAI22S $T=575980 245400 1 180 $X=572260 $Y=245020
X771 748 1 760 148 750 749 2 OAI22S $T=582800 245400 1 180 $X=579080 $Y=245020
X772 164 1 163 162 763 160 2 OAI22S $T=593960 255480 1 180 $X=590240 $Y=255100
X773 164 1 166 162 768 163 2 OAI22S $T=597680 255480 1 180 $X=593960 $Y=255100
X774 164 1 168 162 772 166 2 OAI22S $T=602020 255480 1 180 $X=598300 $Y=255100
X775 748 1 801 183 800 760 2 OAI22S $T=645420 245400 0 180 $X=641700 $Y=239980
X776 184 1 186 183 795 801 2 OAI22S $T=651620 255480 0 180 $X=647900 $Y=250060
X777 802 1 805 187 771 807 2 OAI22S $T=649140 225240 0 0 $X=649140 $Y=224860
X778 802 1 804 187 778 805 2 OAI22S $T=649140 235320 0 0 $X=649140 $Y=234940
X779 189 1 806 187 794 804 2 OAI22S $T=652860 245400 0 180 $X=649140 $Y=239980
X780 189 1 190 187 808 806 2 OAI22S $T=651620 255480 1 0 $X=651620 $Y=250060
X781 813 1 193 194 809 812 2 OAI22S $T=666500 255480 1 180 $X=662780 $Y=255100
X782 812 1 193 194 791 815 2 OAI22S $T=663400 245400 0 0 $X=663400 $Y=245020
X783 197 1 193 194 196 813 2 OAI22S $T=670220 255480 1 180 $X=666500 $Y=255100
X784 193 1 814 194 798 816 2 OAI22S $T=667120 255480 1 0 $X=667120 $Y=250060
X785 828 1 830 831 817 834 2 OAI22S $T=689440 245400 0 0 $X=689440 $Y=245020
X786 846 1 838 844 822 836 2 OAI22S $T=703700 225240 1 180 $X=699980 $Y=224860
X787 845 1 207 845 834 830 2 OAI22S $T=706180 245400 1 180 $X=702460 $Y=245020
X788 845 1 207 212 855 214 2 OAI22S $T=706180 255480 1 0 $X=706180 $Y=250060
X789 853 1 838 853 836 851 2 OAI22S $T=711140 225240 1 180 $X=707420 $Y=224860
X790 853 1 861 853 864 851 2 OAI22S $T=711760 225240 0 0 $X=711760 $Y=224860
X791 863 1 214 859 857 855 2 OAI22S $T=713000 255480 1 0 $X=713000 $Y=250060
X792 861 1 872 868 873 864 2 OAI22S $T=718580 235320 1 0 $X=718580 $Y=229900
X793 918 1 253 918 254 257 2 OAI22S $T=787400 255480 0 0 $X=787400 $Y=255100
X794 1123 1 335 1123 1126 1124 2 OAI22S $T=985180 245400 0 0 $X=985180 $Y=245020
X795 1131 1 1127 1131 1136 1132 2 OAI22S $T=998820 245400 1 180 $X=995100 $Y=245020
X796 1153 1 1154 1155 352 1156 2 OAI22S $T=1017420 235320 1 0 $X=1017420 $Y=229900
X797 364 1 1167 1199 1182 1203 2 OAI22S $T=1040980 245400 0 0 $X=1040980 $Y=245020
X798 1271 1 1252 1278 1276 1281 2 OAI22S $T=1103600 245400 1 0 $X=1103600 $Y=239980
X799 1283 1 1277 1282 1275 1286 2 OAI22S $T=1107320 245400 1 0 $X=1107320 $Y=239980
X800 21 19 22 1 2 474 AO12 $T=256060 255480 1 0 $X=256060 $Y=250060
X801 460 461 28 1 2 486 AO12 $T=263500 235320 1 0 $X=263500 $Y=229900
X802 624 77 80 1 2 638 AO12 $T=409820 255480 0 0 $X=409820 $Y=255100
X803 96 99 650 1 2 658 AO12 $T=444540 235320 0 0 $X=444540 $Y=234940
X804 110 671 661 1 2 679 AO12 $T=471200 245400 1 0 $X=471200 $Y=239980
X805 118 687 690 1 2 119 AO12 $T=487320 255480 1 0 $X=487320 $Y=250060
X806 1031 1029 2 1027 1 1030 AOI12HS $T=874820 245400 1 180 $X=870480 $Y=245020
X807 1045 1047 2 1035 1 1053 AOI12HS $T=886600 255480 1 0 $X=886600 $Y=250060
X808 510 2 512 513 1 AN2B1S $T=298220 225240 0 0 $X=298220 $Y=224860
X809 502 2 512 517 1 AN2B1S $T=301940 235320 0 0 $X=301940 $Y=234940
X810 515 2 512 519 1 AN2B1S $T=303180 245400 1 0 $X=303180 $Y=239980
X811 514 2 512 521 1 AN2B1S $T=305660 225240 0 0 $X=305660 $Y=224860
X812 518 2 512 523 1 AN2B1S $T=305660 235320 0 0 $X=305660 $Y=234940
X813 520 2 512 527 1 AN2B1S $T=308140 245400 0 0 $X=308140 $Y=245020
X814 151 2 748 149 1 AN2B1S $T=567300 255480 0 180 $X=564200 $Y=250060
X815 761 2 802 729 1 AN2B1S $T=647900 225240 1 180 $X=644800 $Y=224860
X816 761 2 193 803 1 AN2B1S $T=663400 245400 1 180 $X=660300 $Y=245020
X817 76 78 1 77 2 620 OAI12HS $T=396800 255480 0 180 $X=393080 $Y=250060
X818 1051 1049 1 1060 2 1059 OAI12HS $T=896520 225240 0 0 $X=896520 $Y=224860
X819 351 1151 1 347 2 1148 OAI12HS $T=1016800 255480 1 180 $X=1013080 $Y=255100
X820 1182 357 1 1178 2 360 OAI12HS $T=1033540 245400 1 180 $X=1029820 $Y=245020
X821 838 835 2 829 207 1 OR3B2S $T=698120 235320 1 180 $X=694400 $Y=234940
X822 7 439 2 1 436 OR2S $T=223200 245400 0 180 $X=220720 $Y=239980
X823 454 8 1 7 440 453 2 MOAI1H $T=242420 235320 1 180 $X=234980 $Y=234940
X824 452 448 449 1 2 454 HA1 $T=243660 245400 0 180 $X=235600 $Y=239980
X825 89 646 647 1 2 651 HA1 $T=428420 245400 1 0 $X=428420 $Y=239980
X826 658 657 665 1 2 670 HA1 $T=455700 225240 0 0 $X=455700 $Y=224860
X827 679 691 698 1 2 701 HA1 $T=491660 245400 1 0 $X=491660 $Y=239980
X828 441 449 442 2 1 XOR2HS $T=234360 245400 0 180 $X=228780 $Y=239980
X829 452 447 456 2 1 XOR2HS $T=238080 235320 1 0 $X=238080 $Y=229900
X830 16 447 459 2 1 XOR2HS $T=242420 235320 0 0 $X=242420 $Y=234940
X831 570 552 576 2 1 XOR2HS $T=342860 255480 1 0 $X=342860 $Y=250060
X832 583 580 587 2 1 XOR2HS $T=351540 225240 0 0 $X=351540 $Y=224860
X833 1097 319 1092 2 1 XOR2HS $T=943020 225240 0 180 $X=937440 $Y=219820
X834 1100 319 1080 2 1 XOR2HS $T=947980 245400 1 180 $X=942400 $Y=245020
X835 1102 319 1083 2 1 XOR2HS $T=949840 235320 1 180 $X=944260 $Y=234940
X836 1103 1101 1094 2 1 XOR2HS $T=950460 225240 1 180 $X=944880 $Y=224860
X837 1104 1101 1084 2 1 XOR2HS $T=954180 235320 0 180 $X=948600 $Y=229900
X838 1061 1046 1062 1 2 1064 MAO222 $T=900240 235320 1 0 $X=900240 $Y=229900
X839 1149 348 1145 1 2 1147 MAO222 $T=1006880 245400 0 0 $X=1006880 $Y=245020
X840 1152 1140 1148 1 2 1135 MAO222 $T=1015560 225240 1 180 $X=1010600 $Y=224860
X841 526 533 541 2 1 525 XOR3 $T=313720 235320 1 0 $X=313720 $Y=229900
X842 666 651 2 655 664 1 656 FA1 $T=462520 245400 0 180 $X=447020 $Y=239980
X843 105 667 2 108 659 1 676 FA1 $T=451980 255480 1 0 $X=451980 $Y=250060
X844 689 669 2 660 681 1 672 FA1 $T=482980 225240 1 180 $X=467480 $Y=224860
X845 683 670 2 675 685 1 696 FA1 $T=478640 235320 0 0 $X=478640 $Y=234940
X846 699 697 2 656 689 1 711 FA1 $T=497860 235320 0 0 $X=497860 $Y=234940
X847 703 709 2 692 701 1 716 FA1 $T=502820 245400 1 0 $X=502820 $Y=239980
X848 708 714 2 700 712 1 723 FA1 $T=509020 245400 0 0 $X=509020 $Y=245020
X849 713 134 2 132 699 1 722 FA1 $T=517700 235320 0 0 $X=517700 $Y=234940
X850 717 724 2 136 713 1 728 FA1 $T=525760 245400 1 0 $X=525760 $Y=239980
X851 720 711 2 730 718 1 734 FA1 $T=530100 235320 1 0 $X=530100 $Y=229900
X852 138 140 2 141 726 1 143 FA1 $T=538780 255480 0 0 $X=538780 $Y=255100
X853 139 721 2 736 733 1 737 FA1 $T=539400 245400 0 0 $X=539400 $Y=245020
X854 731 740 2 742 725 1 754 FA1 $T=548080 225240 1 0 $X=548080 $Y=219820
X855 735 739 2 743 734 1 746 FA1 $T=549320 235320 1 0 $X=549320 $Y=229900
X856 742 750 2 153 715 1 758 FA1 $T=561100 245400 1 0 $X=561100 $Y=239980
X857 152 754 2 759 747 1 756 FA1 $T=566680 225240 0 0 $X=566680 $Y=224860
X858 743 763 2 696 165 1 770 FA1 $T=578460 235320 1 0 $X=578460 $Y=229900
X859 755 751 2 765 767 1 762 FA1 $T=579080 235320 0 0 $X=579080 $Y=234940
X860 764 773 2 775 777 1 169 FA1 $T=590860 255480 1 0 $X=590860 $Y=250060
X861 776 783 2 784 172 1 786 FA1 $T=604500 245400 0 0 $X=604500 $Y=245020
X862 170 785 2 786 171 1 173 FA1 $T=605740 255480 0 0 $X=605740 $Y=255100
X863 773 787 2 788 776 1 175 FA1 $T=608220 255480 1 0 $X=608220 $Y=250060
X864 767 789 2 790 779 1 777 FA1 $T=612560 235320 1 0 $X=612560 $Y=229900
X865 787 178 2 793 797 1 785 FA1 $T=640460 255480 1 180 $X=624960 $Y=255100
X866 789 796 2 795 799 1 788 FA1 $T=647280 235320 0 180 $X=631780 $Y=229900
X867 1017 1026 2 1028 1020 1 1033 FA1 $T=861800 235320 0 0 $X=861800 $Y=234940
X868 1168 1156 1178 1179 2 1181 1 AOI13HS $T=1029200 225240 0 0 $X=1029200 $Y=224860
X869 1176 1206 370 1168 2 1169 1 AOI13HS $T=1045940 245400 0 180 $X=1042220 $Y=239980
X870 1241 1239 387 1161 2 388 1 AOI13HS $T=1072600 255480 1 0 $X=1072600 $Y=250060
X871 60 57 542 582 2 1 MXL2HS $T=354640 255480 0 180 $X=349060 $Y=250060
X872 51 57 564 588 2 1 MXL2HS $T=351540 245400 0 0 $X=351540 $Y=245020
X873 58 57 561 591 2 1 MXL2HS $T=354020 235320 1 0 $X=354020 $Y=229900
X874 61 57 572 593 2 1 MXL2HS $T=355880 245400 1 0 $X=355880 $Y=239980
X875 62 57 568 595 2 1 MXL2HS $T=358360 225240 0 0 $X=358360 $Y=224860
X876 1193 1168 1197 1200 2 1 MXL2HS $T=1039120 225240 1 0 $X=1039120 $Y=219820
X877 447 455 448 445 1 2 HA1P $T=239940 245400 1 180 $X=230640 $Y=245020
X878 15 13 455 11 1 2 HA1P $T=243040 255480 1 180 $X=233740 $Y=255100
X879 1148 1147 1140 2 1 1137 XNR3 $T=1009360 225240 1 180 $X=998200 $Y=224860
X880 592 65 540 1 2 XNR2H $T=358980 225240 1 0 $X=358980 $Y=219820
X881 548 53 2 552 550 1 AOI12H $T=336040 255480 0 180 $X=329840 $Y=250060
X882 573 584 2 580 575 1 AOI12H $T=352780 235320 0 180 $X=346580 $Y=229900
X883 577 580 1 579 592 2 OAI12H $T=349680 225240 1 0 $X=349680 $Y=219820
X884 563 552 1 569 584 2 OAI12HP $T=339760 245400 0 0 $X=339760 $Y=245020
X885 405 2 1 TIE1 $T=1127160 235320 1 0 $X=1127160 $Y=229900
X886 404 2 1 TIE0 $T=1123440 235320 0 180 $X=1121580 $Y=229900
X887 1150 1 2 1158 DELC $T=1019280 245400 0 0 $X=1019280 $Y=245020
X888 849 848 856 847 1 2 215 OA13S $T=707420 255480 0 0 $X=707420 $Y=255100
.ENDS
***************************************
.SUBCKT ICV_34 1 2 3 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 33 34 35 50
** N=69 EP=24 IP=56 FDC=0
X0 11 22 22 1 23 1 2 YA2GSD $T=190720 0 0 0 $X=193570 $Y=0
X1 12 1 1 1 24 3 2 YA2GSD $T=303930 0 0 0 $X=306780 $Y=0
X2 13 3 3 3 25 3 2 YA2GSD $T=417140 0 0 0 $X=419990 $Y=0
X3 14 15 15 15 26 15 2 YA2GSD $T=530350 0 0 0 $X=533200 $Y=0
X4 16 15 10 10 33 10 2 YA2GSD $T=869980 0 0 0 $X=872830 $Y=0
X5 17 10 10 18 34 18 2 YA2GSD $T=983190 0 0 0 $X=986040 $Y=0
X6 19 18 18 18 35 20 21 YA2GSD $T=1096400 0 0 0 $X=1099250 $Y=0
.ENDS
***************************************
.SUBCKT ICV_35
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36 1 2 3 4
** N=5 EP=4 IP=6 FDC=0
X0 1 2 2 2 3 XMD $T=0 1169700 0 270 $X=0 $Y=1109930
.ENDS
***************************************
.SUBCKT ICV_37 1 2 3 4 5 6 7
** N=9 EP=7 IP=12 FDC=0
X0 1 2 2 2 5 XMD $T=0 963780 0 270 $X=0 $Y=904010
X1 3 4 4 4 6 XMD $T=0 1066740 0 270 $X=0 $Y=1006970
.ENDS
***************************************
.SUBCKT ICV_38 2 3 4 6 11
** N=12 EP=5 IP=6 FDC=0
X0 2 3 3 4 6 XMD $T=0 860820 0 270 $X=0 $Y=801050
.ENDS
***************************************
.SUBCKT ICV_39
** N=15 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_40 1 2 3 4 8
** N=9 EP=5 IP=6 FDC=0
X0 1 2 3 3 4 XMD $T=0 449000 0 270 $X=0 $Y=389230
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3 4
** N=5 EP=4 IP=6 FDC=0
X0 1 2 2 2 3 XMD $T=0 346040 0 270 $X=0 $Y=286270
.ENDS
***************************************
.SUBCKT ICV_42 1 2 3 4
** N=5 EP=4 IP=6 FDC=0
X0 2 1 1 1 3 XMD $T=0 243080 0 270 $X=0 $Y=183310
.ENDS
***************************************
.SUBCKT ICV_43
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CHIP out[9] in[7] clk rst_n state[0] state[1] in[0] in[1] in[2] in[3] VCC out[11] GND out[10] out[8] out[7] out[6] out[5] valid resend
+ out[0] out[1] out[2] out[3] out[4] in[11] in[9] in[10] in[8] in[6] in[5] in[4]
** N=3578 EP=32 IP=7384 FDC=0
X0 out[9] 55 729 393 1068 3578 ICV_1 $T=1349740 870270 0 90 $X=1210240 $Y=873120
X1 in[7] 56 2037 3578 ICV_2 $T=0 551960 0 270 $X=0 $Y=492190
X2 3 7 15 18 clk rst_n state[0] 59 state[1] in[0] in[1] in[2] in[3] 2045 57 58 60 67 68 69
+ 70 2038 3578
+ ICV_3 $T=0 0 0 0 $X=139500 $Y=1210660
X3 GND VCC 2038 2092 57 72 2084 73 74 75 2085 78 76 77 79 81 84 82 2086 83
+ 85 80 2087 86 88 87 89 90 3 91 92 2089 97 93 2090 94 95 2096 2098 2093
+ 96 2091 100 101 99 98 103 102 107 2094 104 105 106 2095 59 108 117 109 7 111
+ 2097 2100 2156 115 113 110 114 2099 112 2161 2101 2103 116 2179 2102 2107 2108 2115 2105 2104
+ 124 119 2163 2158 118 120 2162 121 2142 2109 2110 2106 2164 123 2112 2166 125 2111 2114 2113
+ 129 126 2151 2120 2183 174 2116 2182 131 2117 127 168 2185 128 167 2118 2121 2119 2137 187
+ 130 2132 2196 2127 2122 2126 136 2128 122 133 2123 134 2131 2124 2129 135 132 2125 2171 137
+ 138 2165 2175 139 2140 140 157 2130 2184 2138 151 2134 142 2135 145 2136 143 141 147 2143
+ 144 2133 2153 146 2139 158 2148 2157 2172 149 155 2141 2155 148 164 2149 2145 182 153 2144
+ 152 173 2150 156 154 159 2147 2201 160 2167 150 2146 161 2180 2187 162 163 2188 2152 165
+ 166 2154 2173 170 178 169 171 2170 2233 172 175 2218 176 177 2186 2160 2178 2192 180 179
+ 181 183 185 2159 197 184 2209 186 2168 191 188 190 189 2221 2169 213 2174 2200 192 2204
+ 195 194 196 2176 193 214 2177 2190 198 199 2194 2211 2193 200 201 202 2205 244 208 203
+ 204 2229 2195 209 205 2181 2191 206 216 207 2227 211 212 210 215 2223 2197 2199 2198 217
+ 219 220 227 224 218 2207 2202 223 221 2203 2189 2208 226 225 2206 228 2210 229 230 231
+ 232 233 234 2214 236 2216 2215 2217 237 235 239 238 240 242 241 2225 2212 2224 2222 2213
+ 243 2231 245 2228 2230 246 248 247 249 250 251 252 2236 253 2243 2237 256 254 255 259
+ 2234 2239 258 2240 260 2252 257 2242 2244 261 2246 2241 2245 262 265 263 2247 2219 264 2220
+ 2226 2248 273 266 297 268 15 269 278 272 270 271 2257 2254 288 274 275 2253 279 2262
+ 277 276 2258 2259 2260 2256 2263 281 282 283 2266 280 286 285 284 287 2269 2249 2251 291
+ 290 289 292 2271 2304 2274 2268 294 2250 293 267 2235 2278 295 2277 296 2270 2280 300 2279
+ 298 301 299 2281 2283 302 2293 304 2285 2290 2284 303 2287 2286 305 2292 306 307 2276 309
+ 314 308 2267 310 2296 2313 311 2299 2298 312 2300 2301 2303 2275 2305 315 313 316 2294 2232
+ 319 320 321 318 2308 2314 317 2309 2311 2307 2310 322 323 2315 2312 2317 325 324 2316 326
+ 2321 2238 327 2319 328 2330 329 2323 2324 2336 2272 334 332 330 2327 2326 343 333 331 2332
+ 2264 2329 336 2325 335 2255 2088 2333 2291 2331 339 69 2334 341 2341 340 337 344 392 338
+ 2340 2349 2342 2343 347 2345 345 2350 348 346 2348 18 2351 349 350 351 2352 2347 2265 358
+ 352 353 354 2353 360 361 357 355 356 2354 2357 2360 359 2356 362 363 342 364 2335 2361
+ 372 2358 370 365 366 2359 367 2346 2363 368 2365 369 2339 371 2282 2366 375 2364 2362 2322
+ 2368 373 2367 2370 2306 2273 2047 2371 374 2376 2318 2295 2373 2375 378 2372 2302 2385 382 2381
+ 376 2379 377 2380 2383 2382 380 2378 2288 2384 381 2391 2386 2369 2338 2289 2388 384 2389 2390
+ 383 2344 2374 385 2392 2387 2377 386 2355 379 389 2394 2395 387 2337 388 390 2320 2396 2393
+ 2297 2328 391 2397 2045 out[11] 393 2261 3578
+ ICV_6 $T=0 0 0 0 $X=139500 $Y=1086700
X4 GND VCC 71 2084 394 395 397 2398 396 2399 747 2400 2049 2048 398 399 400 2046 402 401
+ 411 2455 404 405 2401 2408 2402 406 2412 408 407 409 2404 2054 410 403 2406 2407 2415 2418
+ 2414 412 2410 2403 413 2411 414 2405 2409 415 2417 416 2413 417 421 2416 420 418 419 2419
+ 2442 422 425 2421 2422 426 2424 2423 428 427 431 57 423 3542 72 2426 429 430 70 432
+ 2425 424 2431 2427 74 2428 2420 73 2429 2435 75 2443 2430 2432 2459 2440 461 439 436 2434
+ 2433 434 435 2437 2469 2438 2436 2439 437 440 438 2446 2468 2085 77 470 76 467 67 78
+ 79 442 2441 80 81 2454 441 2447 68 2086 443 2444 444 2463 2449 445 2452 2453 2445 2456
+ 83 447 2451 2448 84 449 2450 85 448 2484 2464 450 2088 451 86 2087 2457 88 87 452
+ 89 2489 455 2458 453 2465 454 82 477 456 465 482 458 2470 90 459 2460 2474 2461 460
+ 2462 466 91 92 2089 446 464 481 2466 457 2467 2477 95 462 469 2471 93 94 2473 488
+ 2476 471 2480 2090 96 472 97 2091 100 484 98 474 2475 99 2111 475 476 2093 2486 478
+ 2478 479 102 480 2094 103 106 2482 2490 104 105 2095 2499 463 483 108 485 486 101 107
+ 110 114 2485 487 490 2487 2096 2102 2491 2488 2098 2097 2483 111 113 489 112 115 2101 496
+ 494 2107 492 118 117 493 491 2492 2104 2493 119 497 2496 498 495 120 499 501 506 121
+ 500 507 502 122 133 503 2112 123 504 2495 505 124 2494 510 2497 2110 518 126 129 2106
+ 2116 509 2118 512 508 127 511 513 2119 128 2508 515 514 2509 131 132 473 2498 130 134
+ 519 136 516 2479 517 138 2125 521 520 2505 2502 2523 2504 2506 139 2510 2134 522 2129 2503
+ 2517 2516 529 2501 2507 2576 2572 141 524 2570 2138 525 2133 142 526 143 527 2136 144 162
+ 528 2139 2513 145 2512 2143 147 146 2511 530 148 149 2521 2121 2514 151 531 2117 150 2522
+ 154 2147 542 164 152 2144 153 2520 2515 2126 157 155 2146 533 2518 158 2131 532 173 2145
+ 535 160 541 159 536 538 2527 2153 2152 163 2148 161 557 537 546 174 539 2154 534 544
+ 540 165 125 166 181 167 2099 543 2113 168 169 2120 170 171 2500 2156 2157 2158 2100 175
+ 2159 177 548 545 109 182 178 184 2160 2105 2528 468 2050 2542 549 179 2472 2162 185 180
+ 2553 2163 2141 2150 176 550 137 2165 2526 2524 2169 547 551 183 552 2161 553 2530 554 2556
+ 2164 555 2533 559 566 188 2525 2166 2532 116 558 2481 2174 2172 556 190 560 186 561 189
+ 2189 192 2519 2529 2173 193 194 187 195 135 2103 2170 2122 196 2115 2176 2535 563 2171 2177
+ 2114 2181 197 562 2128 2151 199 564 2534 198 2179 2124 2178 214 2167 567 2183 2180 2137 200
+ 565 2108 201 570 568 2195 204 2127 2132 2142 2531 2185 2184 208 2187 572 2536 2182 202 2109
+ 2188 2135 571 2175 203 205 209 2537 172 573 206 574 575 576 578 2538 577 588 569 2540
+ 2186 2190 210 207 579 2539 212 2541 2192 211 2140 2196 581 2123 580 2557 213 216 2223 2543
+ 585 2197 215 2198 222 217 2552 2562 218 219 2545 2199 220 582 2544 583 2546 140 584 2547
+ 2627 221 2548 523 2549 2551 2216 2200 2550 2203 2130 227 2215 587 224 2201 223 231 2193 156
+ 586 2202 2208 226 225 589 2204 2207 590 228 591 2205 230 229 2206 2210 232 2168 2566 595
+ 594 592 593 598 2209 2155 238 2211 234 2194 2213 2149 2212 596 597 2564 243 2560 2214 235
+ 2224 236 233 237 2563 2565 191 2647 599 2219 2575 2217 600 604 2247 602 2225 2220 2226 2567
+ 239 603 2569 2221 2568 605 2571 2222 240 2574 241 606 2573 2228 607 242 610 2580 615 948
+ 608 609 2577 2191 2227 611 245 246 2230 244 252 248 2231 250 612 253 601 2229 613 247
+ 2232 2218 2237 2236 2233 2275 614 2051 2234 2578 254 2582 249 251 617 293 2581 616 2586 2583
+ 2235 2321 618 2319 2579 2585 2558 2555 2601 628 328 2588 2587 619 2591 2584 2554 2612 2600 2606
+ 620 2603 255 625 629 2559 2592 256 621 2593 2590 257 258 2239 2598 259 2238 2561 2243 2240
+ 2594 2589 626 260 622 2241 2599 623 624 2595 2597 2596 2244 2276 627 2242 2250 261 2617 2615
+ 2246 2245 264 2608 2602 2268 262 630 2610 2605 2609 2619 2255 265 631 2604 2611 632 263 2607
+ 267 2614 2251 2249 2613 2264 633 2248 2631 273 634 309 635 2616 266 2625 2620 637 2618 2267
+ 272 268 638 269 2254 2621 2259 270 2624 2253 2252 640 2629 2260 2256 271 2626 2258 2628 275
+ 274 639 2262 276 277 279 2257 641 2263 278 636 281 280 653 2623 2632 2633 642 282 2622
+ 284 2351 2265 2266 283 643 644 2270 286 285 645 2269 287 2278 646 2634 291 288 648 647
+ 2635 2271 289 2311 290 649 2280 295 2630 2274 2636 2272 650 2318 2345 651 652 296 2342 371
+ 294 2273 2364 2326 292 2304 654 659 2384 298 2371 2289 2281 2279 2638 655 2277 2639 300 657
+ 656 2282 2375 658 2283 2383 299 660 297 2640 2292 2290 2651 661 301 302 2325 2642 2288 2286
+ 2284 303 2641 304 2643 2296 662 2285 305 2303 2293 2287 2644 388 2291 2297 2302 2646 2637 668
+ 331 2299 306 2294 308 307 2649 2298 663 2295 2648 2645 315 2300 311 664 665 2650 2301 312
+ 2652 310 677 667 666 313 318 314 670 669 316 2322 317 365 2655 321 671 2305 2306 672
+ 673 2653 2310 320 674 325 2323 2312 2308 2309 345 2656 319 322 2654 675 326 2314 330 323
+ 676 2397 2316 2315 2313 2317 2307 2320 324 2348 678 680 679 2392 332 329 688 682 390 2661
+ 2344 327 2328 333 2324 681 684 387 334 2658 2657 335 336 683 337 2327 2668 342 2662 2681
+ 685 2393 686 338 2390 2330 2660 2332 2666 2331 2334 363 2329 339 2679 2333 2359 356 2336 2665
+ 2341 2335 2659 340 2684 687 693 694 343 341 2338 695 2361 2670 344 2337 2669 689 691 2343
+ 2667 690 2355 2346 692 2672 2339 2349 2340 2674 347 2671 2673 2676 346 2350 2675 2678 2353 350
+ 698 2685 697 2357 2352 696 352 351 359 699 2347 353 2695 366 349 360 354 2366 2354 2677
+ 2368 357 2356 2683 358 355 701 708 361 700 2680 2360 702 2682 2365 703 2363 370 364 367
+ 2053 2358 362 706 704 2362 2367 705 374 707 2370 712 2374 2691 373 2686 372 369 2378 711
+ 348 709 2369 2377 368 386 2395 2372 710 2373 2379 714 2376 382 375 713 2386 385 376 2380
+ 715 716 2381 2689 2047 2382 2694 378 717 379 2687 2385 389 718 2387 2690 381 2391 2688 720
+ 719 380 2394 2389 728 383 2692 377 2396 721 722 2388 7 1067 726 2693 391 384 724 723
+ 2663 725 727 2696 2697 392 729 out[10] 393 2664 3578
+ ICV_18 $T=0 0 0 0 $X=139500 $Y=900220
X5 GND VCC 56 395 733 394 2709 731 397 2398 732 396 2399 734 2701 2049 398 735 2698 2712
+ 730 399 2700 736 2699 737 400 740 2706 401 738 739 742 402 2445 753 2404 403 404 405
+ 2402 409 741 2704 2401 406 407 743 408 2703 744 2403 2410 410 2407 2405 2702 2411 2063 2409
+ 2447 2414 415 411 2408 412 2713 748 2705 746 419 2406 416 417 2711 2415 413 2417 2416 2420
+ 2708 2046 418 2707 749 2413 414 750 2418 751 421 2037 2412 422 420 754 2710 2716 2048 426
+ 423 2419 424 425 2422 2055 2421 755 2424 756 427 428 2714 2425 2400 2427 429 757 430 2426
+ 431 432 433 2429 2428 2431 2433 2432 2430 760 758 441 2434 439 436 434 2715 763 2436 435
+ 2718 759 761 2438 2435 2440 437 752 2469 762 438 3542 2437 470 2719 2439 2826 464 2449 2441
+ 444 2717 765 457 440 2443 2442 442 764 767 2803 2468 443 2837 445 2446 2799 768 766 2444
+ 769 447 770 2448 2720 2452 2825 446 771 2453 448 2451 449 2450 451 450 2454 772 782 2455
+ 453 2728 452 2771 775 774 2723 454 2465 455 2729 780 778 2462 2721 776 2460 2808 2461 456
+ 790 2724 459 460 2463 2811 2471 777 461 773 2725 2464 466 458 2476 462 873 465 463 2467
+ 2726 2722 2459 781 2466 2727 467 779 2470 2730 468 469 2828 2731 472 2472 783 2483 481 784
+ 785 2473 2475 473 786 474 787 2474 488 471 475 2479 2789 476 789 2480 2477 2478 788 477
+ 478 483 479 2500 2733 798 793 792 2481 482 796 812 794 2736 791 802 2732 809 2738 484
+ 2734 486 795 2737 2750 485 2485 2735 487 797 2751 2525 804 2742 2486 800 2488 2754 2530 799
+ 564 2752 801 2740 2487 2519 2755 2739 489 803 493 490 808 2748 492 491 2514 2492 2743 494
+ 495 805 501 496 499 806 2494 2498 2493 497 807 500 2741 810 503 506 498 813 504 814
+ 2496 2744 824 811 2491 509 817 507 823 2502 508 815 502 2746 2747 816 820 510 2749 511
+ 523 819 512 2497 2050 505 821 2490 2548 513 514 825 846 519 822 515 2499 516 525 827
+ 847 2759 517 518 818 826 2756 524 831 521 2783 520 830 2501 2506 526 2505 829 2504 2503
+ 828 832 529 2507 522 2762 833 842 2508 834 527 837 2509 836 2495 528 2512 838 2511 840
+ 531 530 2515 841 839 2520 2513 2767 2510 844 2769 2516 843 2517 532 845 2522 2898 851 945
+ 533 849 540 534 2772 538 536 848 2482 480 2521 850 2778 852 2922 537 539 853 545 535
+ 542 2518 543 854 855 546 544 2523 856 857 2784 548 541 2528 2801 858 2795 859 2802 860
+ 547 2926 861 2780 862 865 864 2776 863 2785 549 867 2781 869 2793 866 2782 868 2909 2524
+ 2790 553 2794 2797 2526 2787 2760 835 2817 870 562 551 552 871 2765 554 876 555 2779 2527
+ 872 2804 556 557 875 2899 559 874 2805 2875 2936 558 560 2529 2809 2788 2536 2806 2812 2851
+ 879 561 563 2821 881 2822 882 877 880 2820 883 889 3549 2815 884 567 2855 886 2768 885
+ 2836 2190 2813 2824 2745 565 571 888 2873 2830 566 887 2532 3547 2773 3545 891 890 2791 2774
+ 3546 2807 2887 2534 892 2835 2533 570 2770 893 569 2800 895 2832 894 2834 2758 896 3552 2757
+ 2823 2539 2766 568 2535 903 897 2814 898 2831 2763 899 572 901 902 905 2537 904 994 575
+ 573 574 2538 576 577 2846 906 2761 578 907 910 913 2764 2552 2557 2540 911 912 2541 908
+ 925 2847 579 2854 2816 581 909 2849 2545 2544 2543 583 915 2857 580 2547 916 2546 914 2549
+ 608 918 582 584 932 951 585 2753 920 2551 2584 587 917 921 922 923 586 2550 919 924
+ 2542 2561 2883 588 927 2860 2554 2864 599 2853 2866 3554 2553 2555 589 930 926 2869 931 1226
+ 2556 594 2559 590 591 2558 2871 2577 929 593 592 937 2874 934 2863 2858 2560 2876 2775 935
+ 2877 2852 2878 900 2810 941 936 2910 2880 938 597 2568 3544 595 940 2792 939 2881 2867 2565
+ 2890 2859 598 2884 947 2563 943 949 2845 600 942 2889 596 2833 2885 1241 2564 602 2861 601
+ 2886 2882 944 2567 2569 2912 2566 2896 2562 603 2585 2796 604 2865 946 2571 2573 2921 2901 3553
+ 607 2872 948 605 2894 2888 2827 950 2574 2842 2913 2798 2891 2777 2572 952 2786 2892 2893 2840
+ 3555 610 609 2575 2576 2570 2895 2580 973 2897 606 953 611 2900 959 2915 2907 612 2908 2902
+ 2903 954 956 2848 2906 955 2905 614 2904 3556 2856 2819 3551 619 957 975 616 958 2956 2868
+ 618 2957 2581 2841 2964 615 2920 2586 2589 878 2604 617 3558 2051 960 3557 3548 2582 2579 2583
+ 2919 2844 613 961 2961 933 620 2591 2870 2578 2862 962 928 2850 2911 2914 629 2916 621 637
+ 3559 2818 626 622 2621 2595 2609 2839 2829 2879 630 625 2600 2843 2056 627 628 623 2602 2838
+ 2592 963 972 964 965 3550 2603 967 2917 2918 2610 631 2928 970 969 632 2624 633 966 2605
+ 2614 2612 968 1014 2616 999 634 635 971 624 638 976 636 2618 2622 974 2966 2632 2923 983
+ 2620 2623 2924 981 640 2625 2619 979 2925 977 2628 639 2627 2927 978 2626 980 2630 2931 646
+ 641 2930 2932 984 645 642 982 648 985 652 653 643 2929 644 986 2940 650 2942 2933 2934
+ 647 987 2634 2935 2939 649 2945 988 2635 2937 2633 2636 993 989 2938 2941 651 991 2949 659
+ 992 2946 2943 2944 990 998 2947 2948 654 655 2639 658 660 657 995 997 656 2951 2950 2952
+ 2640 2644 2954 661 2651 1000 1063 2645 1002 664 2653 1066 662 2955 1011 2648 670 2647 1003 663
+ 1001 666 2649 2953 667 669 668 665 1005 677 1008 1018 671 1013 2650 2962 1006 2652 672 1045
+ 996 2656 673 1007 674 2052 2057 676 1010 675 1009 2959 2655 2960 2654 2958 2967 1004 1012 1016
+ 678 1017 1015 2963 680 679 682 681 1020 2658 1065 683 2661 1019 684 1022 2668 1021 2657 1026
+ 1023 2666 2965 686 685 2970 2981 2663 2670 2980 1024 2660 2669 2968 1028 2659 2696 2662 2671 687
+ 2665 1025 688 690 2672 2679 1027 2684 693 2973 689 2677 1029 2667 2969 691 1030 2673 2674 699
+ 2678 1039 694 1031 695 697 696 2971 2675 2972 1032 1037 1033 692 2683 2686 2676 1034 698 1035
+ 2680 1043 701 2681 2682 2974 2979 704 703 700 1036 1038 2685 1040 702 1042 1048 706 1044 1041
+ 707 1057 1046 1047 2692 705 709 708 1052 1049 1050 2975 2690 2977 2976 712 710 711 1051 1053
+ 1054 1058 1055 713 714 715 720 716 2053 2689 2688 717 1056 718 1059 2694 2687 2978 2693 721
+ 2691 1060 728 2695 727 719 725 722 2697 1061 724 1062 1064 726 723 392 55 3578
+ ICV_23 $T=0 0 0 0 $X=139500 $Y=723820
X6 GND VCC 1069 2982 2983 2984 730 2988 2985 1073 2709 2986 1070 2989 2987 731 733 732 736 2992
+ 1072 2990 734 742 735 1075 1074 2699 1071 2698 737 2700 739 738 740 2991 743 1077 2701 2456
+ 1078 2710 741 2994 1079 2996 2063 745 752 1076 744 750 2702 1080 2704 758 2705 2993 1081 2706
+ 1084 1083 746 1082 2708 747 761 3080 1103 749 748 1085 2997 2058 2054 2995 1086 2999 2703 2037
+ 751 1088 753 2711 754 3000 1091 2068 1089 3082 3004 1090 3001 2712 2713 1087 755 1101 1092 2998
+ 763 2423 2072 3002 3003 2714 1093 756 2715 757 1095 759 1098 1096 1097 2055 2412 3005 2719 2716
+ 3007 1100 2718 3014 3015 3034 2707 760 2720 2717 1094 762 770 1102 764 3033 3006 3020 1105 1104
+ 3019 1107 766 767 768 2721 769 765 3008 1106 1110 3018 2457 1099 772 1108 3021 773 3016 2458
+ 2724 775 1109 3009 1123 3011 778 774 771 1112 2088 3010 776 1954 1111 1114 3012 1113 3071 2726
+ 1118 2722 809 3013 777 1115 3141 2725 779 1116 2723 780 781 1117 787 3017 2728 2730 783 782
+ 3022 1119 786 2729 784 1120 785 2731 1121 3024 3025 788 789 3026 1122 3023 790 1124 1130 3027
+ 1127 796 1125 2734 791 1126 2733 792 2732 1128 793 3028 2736 794 795 799 1142 3030 1129 797
+ 801 798 1131 800 808 1137 1132 2739 802 803 1133 804 2743 2741 1135 805 1136 1134 1140 3031
+ 1138 806 1141 1139 807 3032 2744 1150 810 3035 3029 2727 3036 811 3038 1146 3037 2738 812 1145
+ 813 1147 814 2745 1144 1143 2774 827 815 817 819 2749 818 1148 2060 2746 3039 1149 820 1153
+ 825 1152 822 816 821 1161 3040 2747 823 569 846 3041 2750 824 1154 3042 3043 2531 1155 826
+ 3047 1156 3044 828 2737 1151 919 1157 2740 1158 3056 829 2753 830 2832 3046 1159 1162 2756 2762
+ 2752 2758 831 1163 835 3048 2754 2751 1164 1166 832 2742 2735 2760 2748 1165 2834 2755 833 3049
+ 2759 834 3051 3050 2757 1167 836 1168 3045 2761 838 837 1169 849 1171 2764 1170 1172 2059 1178
+ 2763 839 2772 841 3053 840 2766 2765 1160 842 3052 843 1174 2768 2773 844 2769 1173 3054 2767
+ 2770 3055 2858 914 845 1187 851 847 848 2775 2854 853 1181 2798 1179 2784 2776 1175 850 1176
+ 2777 2778 3057 2833 1177 1189 852 2781 2780 2779 900 2797 2795 855 2885 2782 3058 2787 2786 2793
+ 2863 2791 2810 2816 2783 854 3059 2788 2840 2794 2785 860 908 3544 2847 2800 952 1186 857 862
+ 858 3060 2790 2807 2857 856 1180 2892 859 2906 3061 861 1194 1198 1182 3545 866 3062 2856 2792
+ 1183 864 1184 865 2796 867 863 1185 2845 3551 868 869 3064 2842 870 1191 1188 3558 871 2844
+ 906 3063 2823 3065 1190 2789 2841 872 3548 2849 3546 3066 2802 941 2824 2799 2801 2803 2862 2870
+ 2808 961 2804 2881 2813 899 1192 2822 2806 1193 873 3557 2848 2850 2811 2839 1197 879 2809 874
+ 2821 2021 2805 876 3556 2056 2814 875 1561 881 2818 1195 3072 882 2865 2815 2812 877 1196 3547
+ 2829 2843 3067 878 3068 3553 3549 1203 2875 2819 2827 912 880 1199 2853 3550 2820 2911 3555 883
+ 2868 2846 884 1230 2866 2852 2484 894 3070 885 1229 3074 2637 2867 2826 2771 2825 2828 924 2489
+ 1200 886 888 1201 2831 1210 889 2830 1202 1204 891 892 2872 2836 3552 890 3073 893 1549 898
+ 887 2835 895 1205 2838 2817 2837 896 1214 897 2861 3088 1234 2918 2859 3076 1206 1207 902 903
+ 1208 911 3086 905 1209 1211 904 60 3085 994 3079 3075 907 909 910 2851 1212 2855 913 1213
+ 1216 1215 916 901 1217 915 1218 2902 3078 918 917 1219 1220 931 2860 926 921 922 3081 1225
+ 3083 920 923 1223 3094 2864 925 1221 927 1222 2916 1224 3084 932 930 929 928 3087 3090 2092
+ 1231 3089 2873 1227 3093 935 1228 3091 934 933 940 938 936 2879 1235 937 1232 2882 939 946
+ 1240 942 2883 2890 1233 3554 943 944 1236 1239 2914 1247 609 2562 2896 3095 1237 1238 2880 950
+ 3559 3105 3100 3099 2570 1241 1255 3104 945 1242 1250 2889 3098 947 1243 3097 2576 3096 948 2887
+ 2888 2574 951 2891 2925 2893 1244 1246 2931 2895 949 3101 1245 1248 2897 1249 953 2901 2899 956
+ 3103 2904 2900 954 3102 2908 960 955 2903 2905 2907 957 3110 958 1251 989 1252 1253 3108 1254
+ 1257 3107 2910 2913 959 1015 964 3111 1256 2917 1258 3117 3109 3116 3113 2951 3112 1259 982 3106
+ 3114 3123 2588 2598 1261 3069 1262 1260 2587 966 2594 968 969 1264 2599 970 2928 2606 3120 2593
+ 2607 2611 2920 2590 2597 2613 1267 1263 967 2601 2919 1265 971 3115 2617 2615 3119 2922 973 1268
+ 2608 3121 3126 2596 1266 1270 975 3125 1269 1272 976 974 3124 3118 3122 2924 977 2909 1275 2915
+ 3133 1273 1277 2926 3127 3128 979 1274 3077 3134 3130 3131 2629 972 3129 1276 3135 1279 981 2923
+ 1278 980 3132 1280 2929 2631 1286 985 3092 3163 984 1281 3136 983 1282 963 3137 2932 1284 1285
+ 987 1290 986 3139 3138 2933 3142 3140 2937 2936 1287 1288 2943 1289 2941 990 2947 995 988 991
+ 993 992 1292 1291 1644 2945 3145 3146 3143 3192 2948 996 1293 2061 3158 2949 3144 2057 1294 965
+ 1000 1295 2638 997 3147 1296 1297 2953 1310 2954 3159 1298 1556 1326 998 2641 2643 3148 3182 2642
+ 2646 3162 1002 1001 3184 3149 3151 1557 1299 3150 1301 2955 1300 1003 1302 1004 1005 1304 1305 1303
+ 3155 1312 2062 1306 3170 3153 3154 1006 1307 3152 3156 2958 1308 1009 1007 2959 1008 1309 3157 3160
+ 1010 3179 2960 1011 3172 1311 999 1314 1013 1012 962 1014 1315 3165 1715 2961 1016 2957 3161 3207
+ 1316 1317 1018 1017 2963 2967 683 2964 1319 1318 3166 3178 2956 3167 2971 1322 2962 1019 1325 2965
+ 3169 1313 3183 3199 3168 1020 3175 3176 3189 3206 1320 3173 2966 1321 1021 3174 3171 1022 1323 3181
+ 1027 3180 1324 1023 1024 2968 3187 3186 3188 3185 1328 1327 1026 3193 1329 3177 1339 2973 1330 1029
+ 3190 2969 1331 1028 1687 3164 1035 1030 1332 1333 2972 3191 3196 1031 1033 1032 1334 1038 1034 3194
+ 3197 1036 3195 1335 1037 1337 3203 1336 1338 1039 3198 1042 3202 1040 2978 3208 1041 1043 1045 1344
+ 2975 1044 1342 2974 1048 1343 3200 1046 2977 1341 1340 1050 1049 3205 1053 1052 3201 1051 1047 1347
+ 1054 1059 1345 1346 1349 1055 1056 1350 1060 1348 1058 1352 1353 1356 1064 2976 1351 3204 1354 1358
+ 1061 3210 1062 2979 1063 1065 1066 2981 2980 1355 2970 out[8] 1357 393 3209 3578
+ ICV_29 $T=0 0 0 0 $X=139500 $Y=533370
X7 GND VCC 56 3211 3212 2989 1069 1359 2988 2991 1362 2984 2985 1073 1360 2982 1361 2983 1074 1070
+ 3214 1071 2986 3213 2990 1364 1363 1365 2987 1072 3215 1370 1366 1367 1372 1369 1368 2058 1075 1076
+ 1375 1371 2994 1077 2992 1378 1078 3216 1079 2995 1081 2993 1374 1376 1377 1080 1082 1379 3217 2996
+ 1381 1382 1084 2997 1083 1383 1380 3218 1385 1085 1384 1386 1387 1388 1092 2998 1390 1389 1090 1087
+ 1086 1373 2999 1391 1089 3000 3001 1088 3002 1091 1392 1393 3003 1093 1394 1395 1396 1397 1094 1095
+ 1096 1097 1098 1099 1398 3219 3237 3236 1101 1100 1399 1400 1102 1720 1103 3007 1416 1401 1104 1109
+ 1106 1402 1105 1403 3227 1404 1107 1406 1405 1407 1439 1108 1408 1409 765 1410 1411 1110 3222 1412
+ 1111 3009 3223 1418 3224 1413 1414 1112 1415 3221 3226 3006 3225 3014 1417 1419 1113 1114 3008 1115
+ 3013 3018 1116 1421 1422 3017 3015 1117 1118 1423 3233 1119 3019 1428 1424 1437 1120 1425 3229 3016
+ 3020 3230 1430 1126 1426 1433 1427 3023 1420 1121 1429 3021 1752 3022 1431 3231 3026 1432 3024 1122
+ 3232 3025 1124 1123 1434 1435 1436 3027 1438 3028 1125 1127 1510 1128 1440 3234 1441 3238 1129 1442
+ 1130 1444 3240 1443 3239 3029 1445 3030 3242 3241 3053 3245 1447 1451 1453 1131 1446 1132 3220 3244
+ 1449 1448 1133 3246 1136 1142 3235 1450 1137 1134 1458 1135 3033 1452 1139 1140 1454 3031 3032 2074
+ 1141 1455 3247 1459 1138 1456 1457 3036 3035 3251 3037 3249 1460 1147 1498 1150 1790 1148 3039 1461
+ 816 3038 1143 1464 3228 1146 1144 1145 3248 3250 1462 1463 1465 1466 1160 1151 3041 1152 3040 3043
+ 3252 1153 1156 3049 3045 1467 3253 1154 1798 1469 1470 1163 3056 1468 3042 1471 1149 1155 1472 1473
+ 3044 3046 3254 1157 1158 1159 2060 1161 3256 1164 1474 1475 3047 1476 1165 1166 3048 1162 3262 1490
+ 3258 1477 1478 1480 3257 1178 1169 3050 1171 3260 1172 3265 1167 3259 3275 3051 1168 3285 3276 3264
+ 1481 3294 2059 3052 1170 3280 3261 1479 3267 3263 1496 3054 1482 3059 3266 3268 1484 3269 1485 1486
+ 1487 1488 3270 1489 3271 1173 1174 3055 1491 1492 1176 1493 3273 1499 3255 1494 3272 1495 3274 1175
+ 3057 1177 1187 1497 3064 1179 3058 3277 3278 1501 3279 1500 3063 3282 3281 3060 3284 1504 1502 3283
+ 1180 3286 1194 1181 1182 1505 1506 3062 1507 3068 1508 1183 1188 3289 1509 1184 3061 1185 1511 1503
+ 1513 3243 3288 1196 3287 1514 1186 1512 1189 3067 1515 3290 3065 1190 1191 1192 1516 1193 1518 1519
+ 1517 3291 1197 1195 3066 3292 1520 3293 1198 1199 1265 3305 1524 1522 1521 1200 3069 3115 1201 1203
+ 1202 3296 3295 3106 1528 1204 1525 1526 1527 1529 1228 3297 1530 3302 1531 1205 3301 1532 1206 3299
+ 1207 3298 3300 1208 3310 1209 3122 1534 3304 3307 1540 1537 1214 3303 1210 3118 3073 3072 1535 1211
+ 1538 3132 1212 1536 1545 1266 3306 3311 1215 3092 1216 1543 1541 3077 1218 1213 3308 1542 3309 1539
+ 3312 1533 1544 1219 3078 1523 1220 3084 1227 1222 1546 1225 1223 3081 3089 3083 3090 1221 2869 1226
+ 1548 1547 1217 3094 1224 3087 2871 2874 3091 1229 1230 1552 2876 3093 1578 1232 2878 1231 1551 2877
+ 1550 1237 1554 1233 1236 1234 1239 2884 1235 2886 1555 1238 3313 1553 1247 1558 1559 3095 1240 3314
+ 3317 3097 1560 1242 3100 3096 1241 1562 3099 3315 1243 3105 1244 1249 1572 2898 3316 1579 3098 1245
+ 1564 2894 3318 3101 1246 1248 1565 1584 1254 1567 1568 3103 3319 3102 1250 3112 1566 3320 1563 1570
+ 1569 1571 1251 3108 3107 1252 1573 3109 3321 1574 3111 3110 1257 1255 1253 3322 1256 1575 1258 1576
+ 1581 1259 3113 3325 1580 3326 3324 3333 3329 3114 1260 1577 3335 3328 3323 3334 3327 3330 1261 3104
+ 3331 3332 3336 1583 1262 3116 1588 3117 1585 1590 1263 1586 1589 2912 1587 3120 1591 1267 3337 1596
+ 3121 3339 1268 3139 3123 1594 3342 1270 1271 1272 1269 1597 3341 1595 1592 1593 3340 3358 2921 3343
+ 1264 1287 1273 3344 3124 3347 2064 1598 1599 1274 3126 1275 3338 3346 3128 3127 1601 1600 3345 1279
+ 1277 1607 1276 1278 1611 2927 1603 1292 1606 3131 978 3119 1605 1608 3350 3125 3129 1280 3135 3349
+ 1609 2061 3130 1610 3134 3133 1604 1281 1620 2930 3359 1612 1285 3352 3136 3137 3138 3356 1284 1282
+ 3351 1283 1615 1614 3354 1286 1613 1617 2934 1295 3355 2940 1619 1616 1602 1289 1621 2938 2935 3357
+ 2939 3353 3140 1618 2942 1290 1288 1622 1623 2946 3376 1637 2944 3360 3348 2065 1624 3362 3369 1310
+ 3147 1294 3361 1625 3145 1631 1626 2952 2950 3151 1627 1296 1628 3364 3368 1629 1297 1630 3363 3366
+ 3367 1298 3365 3382 1632 3402 1633 3371 1299 1636 1655 1640 3374 1634 3384 3378 3150 3385 1638 3149
+ 1639 3383 3370 3161 1641 3377 1642 1635 3373 3379 1305 3407 1304 1301 3375 1643 1646 3386 1645 1303
+ 3392 1300 1647 1651 3401 3390 1688 1648 3381 3399 3380 3398 1653 1302 1649 3387 1650 3400 1652 3389
+ 3388 1658 1654 1662 3396 3391 3393 3394 1657 3397 3428 3395 3408 1306 3403 3404 1656 1307 3155 3406
+ 1308 1660 3405 3156 3153 3417 3416 3158 1311 3411 1321 1314 3409 3144 3420 1668 3425 1661 3160 3424
+ 1313 1664 3172 1315 1659 3415 1665 3430 3412 1663 3162 3410 3414 3413 3164 3165 3178 3173 1666 1667
+ 3167 3166 3418 1317 3191 3423 1318 3561 3169 3163 3427 3421 1319 3419 3168 3431 1316 3180 3171 1676
+ 3176 1322 3426 3174 3170 3175 3422 1324 1670 1323 1669 3179 3159 3148 3188 1671 1675 3429 3182 1325
+ 1679 3177 1672 1326 3185 3435 3187 3434 3186 1673 3440 1674 3432 1327 1328 3189 3436 3447 3442 3433
+ 3184 3181 3190 1330 1678 3562 1677 1680 1331 1682 3183 3438 3437 3448 1329 1681 1332 3439 3449 3146
+ 1683 1704 3441 1333 1684 3445 3444 3192 3443 1686 3450 1685 2066 3194 1335 1689 1334 3195 1703 3446
+ 1710 1691 1696 3451 1338 3197 1336 1337 1692 1693 1695 3454 3452 1690 3453 1351 1339 1699 3455 1343
+ 1340 3457 1697 1711 1341 1698 1694 1700 3456 1702 1342 1701 1346 1705 3467 3201 1344 3465 1706 1347
+ 1707 3204 3202 3203 1708 1345 3460 1709 3458 3459 3461 1348 1349 1352 3464 1350 3463 1712 1716 1713
+ 1354 3466 3462 1355 3468 1714 3200 3152 3205 1358 1353 1067 3154 1357 1717 3210 1356 out[7] 393 3372
+ 3578
+ ICV_31 $T=0 0 0 0 $X=139500 $Y=365980
X8 GND VCC 1719 28 3212 1718 1362 1720 1722 1721 1359 3211 1360 1361 1363 1070 1401 1723 1365 1364
+ 1728 1726 1724 1727 3213 1725 1733 1366 3469 1367 3214 1368 1369 1729 1370 1730 3215 3470 1372 1371
+ 3473 3472 1731 1373 1375 1732 1374 3471 1734 3216 1736 1735 3474 1378 1376 1377 1738 1743 1380 3217
+ 1739 1381 1740 2073 1379 1742 1383 3475 1741 1382 3476 1385 1384 1737 1386 1388 1744 1747 1387 1745
+ 1389 1390 3218 1392 1391 1746 1395 1403 1748 1394 1396 1749 1393 1397 1750 1751 3219 1398 1399 1400
+ 1753 1754 1404 1402 1774 1755 1405 1756 1757 1408 1406 3477 3220 1410 3228 1409 2067 1411 3222 1759
+ 1758 3221 1407 1412 3478 3224 1413 3223 1414 1760 3225 1415 3010 3248 3226 1416 3234 3011 1417 3236
+ 1761 1419 1418 3227 1510 1762 1420 1763 1421 1422 1438 1423 1764 1765 3479 1424 3480 1766 1767 1428
+ 3481 1425 3229 3230 1432 3233 1768 1770 1426 3482 3232 1429 3483 1769 1433 3231 1430 2068 1427 1431
+ 1771 1772 1435 1437 3025 1773 1436 1434 1775 1776 1777 3256 1780 1439 3242 1442 3238 1440 3239 1445
+ 1441 1778 1449 3484 1443 1779 3485 3241 3240 1444 3237 3486 1446 1781 3487 1452 3254 3244 1447 3243
+ 1782 1448 3245 1784 3488 1785 3247 1783 1786 1451 1454 3246 1450 1453 1789 1791 3489 1455 1788 1456
+ 1793 1792 1790 1457 3249 1459 1458 1460 1794 1795 3490 1461 1465 1796 1462 1799 1463 1798 3250 1464
+ 1797 1466 1467 1787 3255 3251 1468 3252 3253 1800 1470 1471 1469 1830 1472 1802 1803 1804 3293 3053
+ 1805 1807 1806 3277 3493 1473 1808 3257 1477 1478 1810 3497 3258 1811 1833 3261 1494 1812 1479 1474
+ 1480 1813 1475 1481 3264 3263 1482 1483 1476 3262 3266 3267 1484 3269 3268 3259 1486 3271 1487 1488
+ 1815 3260 1489 1490 3270 1817 1816 1821 1491 1492 3265 1814 3491 1493 3272 1485 1495 1819 1818 3492
+ 3274 3273 1496 1822 1497 1498 3275 1809 1499 3278 1824 3496 1823 2075 3276 1500 1829 3281 1825 3494
+ 3495 1820 1504 3283 1501 3282 1502 1508 3279 1826 1503 1827 3280 1505 1506 1828 1507 1851 1831 1801
+ 3290 3498 3286 3285 3287 3499 3288 3297 1832 3289 2025 1512 1513 1514 1515 3500 1835 1509 3501 1836
+ 1837 3298 1516 3284 1838 1834 1517 1518 1519 1840 1839 1844 3292 1845 3291 1841 1520 1843 1842 1522
+ 3296 3294 1524 1846 1521 1523 3305 3295 1528 1847 1525 1526 1848 3301 1532 1530 1849 1529 1527 3300
+ 1531 3308 1850 1852 3302 1542 1856 3502 1544 3310 1854 3299 1853 1855 3503 3303 1857 3504 1533 3304
+ 1535 3307 3306 1534 1859 1858 1538 1536 1537 1545 1539 1860 1541 1861 1540 3309 1543 3311 1863 3312
+ 1862 3505 1864 1546 1865 1548 1867 1868 3075 2020 1875 1547 58 1869 3088 3506 3079 1549 1870 1871
+ 3076 1866 2069 1550 2022 1873 1874 1552 1879 3313 1872 3074 1877 1553 1554 3071 1551 3086 1880 1555
+ 1876 1558 1881 1882 1556 1878 1888 1557 1559 1560 1883 3085 1884 1885 1561 1562 1886 3314 3070 1563
+ 3315 1887 1564 1897 3316 1569 1891 1566 1889 1892 1890 3317 3318 1565 1893 1567 1584 1579 1571 1895
+ 1894 3319 1896 1568 1898 3507 1899 1570 1572 3320 1900 1901 3321 3508 1573 1903 3004 1576 3322 1574
+ 3082 1575 1905 3509 1580 1906 1577 3323 1578 3510 1910 1908 1909 3326 3327 1907 1581 3511 3324 1582
+ 1911 3328 3372 2055 3325 1904 3512 1583 1912 3329 1913 3331 3513 2714 3330 3334 1585 1914 1917 1587
+ 1915 3332 3333 3514 3336 1916 3209 1588 3515 3335 1918 3080 1586 1919 1591 1589 3413 3516 1592 1590
+ 1068 3345 2707 1593 1920 1922 3337 1921 1902 3338 3517 1594 1923 2031 1596 3339 1925 1595 1983 3518
+ 1597 1924 1598 3342 1600 3519 3343 2664 3358 3341 3352 1927 3340 2716 1928 3344 3347 2261 1604 1601
+ 1606 2033 3349 3346 3520 1929 1602 1603 2034 1599 1930 1605 3348 1607 1932 3350 1609 1926 1612 3354
+ 1931 1610 3034 1608 1933 1934 3351 1611 1935 1622 3012 1936 3521 1614 1613 3353 1939 3522 1937 1938
+ 1616 1954 3355 1615 1617 3357 1618 1940 3005 1621 1941 1620 1942 3359 1943 3356 1626 1638 1944 1623
+ 1945 3141 1624 1946 3360 1625 2065 3362 3361 1641 1627 1949 3365 1628 1950 3364 3367 1636 1629 3363
+ 1947 3366 3368 1648 1630 1948 1631 1639 1633 3369 1653 1634 1951 1968 1632 1635 1953 3373 1952 3370
+ 3382 1637 3375 1640 3371 1646 1642 3376 1293 1645 1957 1955 1643 1644 1647 3379 1956 3374 3380 3378
+ 3402 3523 1974 1961 3383 3395 3391 1651 3384 3385 3388 1958 3381 1652 1650 1959 1963 3386 3401 1655
+ 1649 1656 1960 3377 3399 3393 3397 3394 3400 1283 3389 1658 1962 3403 3387 3142 3398 1965 1657 3526
+ 3406 3396 3392 3405 1964 3524 1654 3404 3390 3409 1671 1966 1662 1663 1660 1291 3415 1661 1664 3407
+ 3143 2070 1969 1659 3414 3412 3408 1665 3417 3416 1666 3419 1970 3411 3410 3180 3525 3423 1967 3418
+ 1669 1971 3424 1312 1667 3422 1668 1972 3421 3425 1309 1976 1973 3426 1673 1670 3427 1678 1975 3561
+ 1672 1679 3433 1977 3538 1978 3429 3420 1674 1979 1980 3430 1676 3434 1981 1677 3431 3432 3436 3435
+ 1675 1982 3562 3193 1682 3442 1680 3527 1984 1681 3528 1988 1986 1987 3440 3438 1684 1985 3536 3441
+ 1989 3529 1689 1990 3444 3439 2066 1683 3530 3437 1711 1685 3449 2082 3445 1686 1687 3531 3447 1688
+ 3537 3532 1991 3533 1999 3450 3448 1691 1690 3534 3446 1993 3428 3196 1992 3443 3455 3453 3454 1995
+ 3452 1692 1994 1696 1694 1996 3451 1693 1998 1997 3535 1697 2000 1695 2001 1700 1699 3456 2002 2003
+ 1698 2071 2004 1710 1701 1702 2005 2007 2006 1705 1704 3467 1703 3457 1706 3458 2010 1707 2008 3464
+ 1708 2009 3459 2011 3462 3460 3539 1709 2012 2013 3461 1712 3463 2014 3465 2015 1323 3540 3466 2016
+ 2017 3199 2018 2062 3208 1714 3157 1318 3198 1715 1716 3206 3207 3468 1717 2019 out[6] 393 3578
+ ICV_32 $T=0 0 0 0 $X=139500 $Y=260100
X9 GND VCC 29 28 1719 1720 1721 1718 1722 1723 1724 1725 1726 1727 1728 1729 3473 3470 1731 1742
+ 1733 3471 1732 3472 1734 1730 3469 1735 1736 1737 3474 1738 1741 1740 1739 2073 1744 1743 3475 3476
+ 1745 1746 1747 1748 1750 1749 1751 1752 1753 1754 1758 31 1755 30 1756 1757 1760 3477 1759 3478
+ 3225 3234 2067 1761 3235 1762 1763 1764 3479 1768 1765 3481 3480 3483 1766 1767 1774 1772 3482 1769
+ 1770 1773 1771 2068 1776 1775 1778 1779 1781 1780 3485 3486 1783 1782 1777 1784 1785 3488 3489 1786
+ 2074 2023 3484 1789 1787 3487 1790 1792 1791 1788 1793 1794 1795 1797 1796 1799 1798 1800 1801 1804
+ 1803 1807 1802 1808 3490 1810 1805 1809 1811 1812 1822 1813 1806 1818 1814 1827 1815 1816 1817 1819
+ 1826 1820 1821 3491 3492 1828 3493 3498 1823 1824 3495 3494 1825 3496 1829 1850 1831 3497 3499 1833
+ 1832 1837 1834 3500 3502 1835 1836 1838 3501 1841 1839 1840 1844 1843 1845 1846 2075 1848 1847 1830
+ 2025 1849 1851 1853 1852 1855 1842 3503 1854 1856 1857 1861 1858 1859 1860 3504 3312 1862 1864 1863
+ 1865 1866 1867 2069 1869 1868 1870 3505 1871 3506 1872 1873 1874 1875 1876 1877 1878 1879 1881 1880
+ 1884 1890 1886 1882 1885 1887 1888 1889 1916 3510 1891 3516 1892 1893 1894 3507 1895 1896 1897 1898
+ 1901 1900 1902 1903 1899 1904 1908 1906 1905 1907 1914 1909 3509 3508 1910 3511 1911 1912 3512 1913
+ 1917 3515 3514 1918 1919 3519 1920 1922 1921 1923 3517 1929 3513 1924 1925 3518 1926 1927 1938 3521
+ 1928 1930 1931 1932 1933 1934 1935 1936 1915 3522 1937 1940 1939 1941 38 1943 1942 1944 1946 1945
+ 1983 1947 1948 3005 1949 1950 1952 1953 1951 3012 1954 1955 1957 3523 1959 1956 1958 1960 1962 1961
+ 1963 1964 1966 1967 1968 3526 1965 1969 2070 3524 1970 3525 1971 1972 1973 1975 1974 2032 1976 1977
+ 1978 1979 1981 1980 1982 1996 1988 3530 1984 1987 1985 1986 3528 1989 3529 1990 3532 3533 1999 3527
+ 2082 3531 1991 3534 1992 2001 1993 1994 1995 3535 1997 3536 1998 2000 2007 2002 2003 2071 3537 2004
+ 2005 2006 2008 3538 2010 2009 2011 3539 2013 2012 2016 2015 2014 2018 2017 3540 1067 2035 393 2019
+ out[5] 3520 3578
+ ICV_33 $T=0 0 0 0 $X=139500 $Y=139500
X10 29 30 31 38 valid resend out[0] out[1] 2023 out[2] out[3] 2032 out[4] 1067 2035 28 2020 2021 2022 1883
+ 2031 2033 2034 3578
+ ICV_34 $T=0 0 0 0 $X=139500 $Y=-56920
X12 in[11] 71 2046 3578 ICV_36 $T=0 0 0 0 $X=-56920 $Y=1087500
X13 in[9] 394 in[10] 71 2048 747 3578 ICV_37 $T=0 0 0 0 $X=-56920 $Y=901000
X14 in[8] 394 56 2054 3578 ICV_38 $T=0 0 0 0 $X=-56920 $Y=724600
X16 in[6] 56 1359 2063 3578 ICV_40 $T=0 0 0 0 $X=-56920 $Y=366000
X17 in[5] 1359 744 3578 ICV_41 $T=0 0 0 0 $X=-56920 $Y=260100
X18 28 in[4] 2072 3578 ICV_42 $T=0 0 0 0 $X=-56920 $Y=139500
.ENDS
***************************************
