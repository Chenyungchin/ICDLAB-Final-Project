module Sobol(
    input         clk,
    input         rst_n, 
    input         start,
    output reg [31:0] res0,
    output reg [31:0] res1,
    output reg [31:0] res2,
    output reg [31:0] res3
);


// ================== reg and wire ======================
reg   [31:0] DVA [0:31];
// reg   [31:0] res0, res1, res2, res3;
wire  [31:0] res0_w, res1_w, res2_w, res3_w;

reg   [31:0] counter;
reg   [4:0] LSZ;

integer i;

// ================== wire assignments ==================
assign res0_w = res3 ^ DVA[0];
assign res1_w = res0_w ^ DVA[1];
assign res2_w = res1_w ^ DVA[0];
assign res3_w = res2_w ^ DVA[LSZ + 2];

// ================== Combinational =====================
always @(*) begin
    for (i=0; i < 32; i = i+1) begin
        if (counter[31 - i] == 0) LSZ = 31 - i;
    end
end


// ================== sequential ========================
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        res0    <= 32'b0;
        res1    <= 32'b0;
        res2    <= 32'b0;
        res3    <= 32'b0;
        counter <= 32'b0;
        // DVA
        DVA[0]    <= 32'b10000000000000000000000000000000;
        DVA[1]    <= 32'b11000000000000000000000000000000;
        DVA[2]    <= 32'b00100000000000000000000000000000;
        DVA[3]    <= 32'b11110000000000000000000000000000;
        DVA[4]    <= 32'b10101000000000000000000000000000;
        DVA[5]    <= 32'b00110100000000000000000000000000;
        DVA[6]    <= 32'b11010110000000000000000000000000;
        DVA[7]    <= 32'b01001001000000000000000000000000;
        DVA[8]    <= 32'b11001011100000000000000000000000;
        DVA[9]    <= 32'b01100101010000000000000000000000;
        DVA[10]   <= 32'b00110010111000000000000000000000;
        DVA[11]   <= 32'b00011001100100000000000000000000;
        DVA[12]   <= 32'b00001100000110000000000000000000;
        DVA[13]   <= 32'b00000110011011000000000000000000;
        DVA[14]   <= 32'b00000011111110100000000000000000;
        DVA[15]   <= 32'b00000001110111110000000000000000;
        DVA[16]   <= 32'b00000000000000001000000000000000;
        DVA[17]   <= 32'b00000000000000001100000000000000;
        DVA[18]   <= 32'b00000000000000000010000000000000;
        DVA[19]   <= 32'b00000000000000001111000000000000;
        DVA[20]   <= 32'b00000000000000001010100000000000;
        DVA[21]   <= 32'b00000000000000000011010000000000;
        DVA[22]   <= 32'b00000000000000001101011000000000;
        DVA[23]   <= 32'b00000000000000000100100100000000;
        DVA[24]   <= 32'b00000000000000001100101110000000;
        DVA[25]   <= 32'b00000000000000000110010101000000;
        DVA[26]   <= 32'b00000000000000000011001011100000;
        DVA[27]   <= 32'b00000000000000000001100110010000;
        DVA[28]   <= 32'b00000000000000000000110000011000;
        DVA[29]   <= 32'b00000000000000000000011001101100;
        DVA[30]   <= 32'b00000000000000000000001111111010;
        DVA[31]   <= 32'b00000000000000000000000111011111;
    end
    else begin
        if (start) begin
            res0    <= res0_w;
            res1    <= res1_w;
            res2    <= res2_w;
            res3    <= res3_w;
            counter <= counter + 32'b1;
        end
        else begin
            res0    <= 32'b0;
            res1    <= 32'b0;
            res2    <= 32'b0;
            res3    <= 32'b0;
            counter <= 32'b0;
        end
    end
end

endmodule